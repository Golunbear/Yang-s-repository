//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2025 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = efx_csi2_tx
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Thu Jun  5 09:44:30 2025
// ***************************************************************************************

`define IP_UUID _csi2tx250605
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)
`timescale 1 ns / 1 ps
module efx_csi2_tx #(
    parameter tLPX_NS = 50,
    parameter tINIT_NS = 100000,
    parameter tINIT_SKEWCAL_NS = 100000,
    parameter tLP_EXIT_NS = 100,
    parameter tCLK_ZERO_NS = 262,
    parameter tCLK_TRAIL_NS = 60,
    parameter tCLK_POST_NS = 60,
    parameter tCLK_PRE_NS = 10,
    parameter tCLK_PREPARE_NS = 38,
    parameter tHS_PREPARE_NS = 40,
    parameter tWAKEUP_NS = 1000,
    parameter tHS_EXIT_NS = 100,
    parameter tHS_ZERO_NS = 105,
    parameter tHS_TRAIL_NS = 60,
    parameter NUM_DATA_LANE = 4,
    parameter HS_BYTECLK_MHZ = 187,
    parameter CLOCK_FREQ_MHZ = 100,
    parameter DPHY_CLOCK_MODE = "Continuous", 
    parameter PACK_TYPE = 4'b1111,
    parameter PIXEL_FIFO_DEPTH = 2048,  
    parameter ENABLE_VCX = 0,
    parameter FRAME_MODE = "GENERIC",    
    parameter ASYNC_STAGE = 2
)(
    input logic           reset_n,
    input logic           clk,				
    input logic           reset_byte_HS_n,
    input logic           clk_byte_HS,
    input logic           reset_pixel_n,
    input logic           clk_pixel,
	output logic          Tx_LP_CLK_P,
	output logic          Tx_LP_CLK_P_OE,
	output logic          Tx_LP_CLK_N,
	output logic          Tx_LP_CLK_N_OE,
	output logic [7:0]    Tx_HS_C,
	output logic          Tx_HS_enable_C,
    output logic [NUM_DATA_LANE-1:0]         Tx_LP_D_P,
    output logic [NUM_DATA_LANE-1:0]         Tx_LP_D_P_OE,
	output logic [NUM_DATA_LANE-1:0]         Tx_LP_D_N,
    output logic [NUM_DATA_LANE-1:0]         Tx_LP_D_N_OE,
	output logic [7:0]                       Tx_HS_D_0,
	output logic [7:0]                       Tx_HS_D_1,
	output logic [7:0]                       Tx_HS_D_2,
	output logic [7:0]                       Tx_HS_D_3,
	output logic [7:0]                       Tx_HS_D_4,
	output logic [7:0]                       Tx_HS_D_5,
	output logic [7:0]                       Tx_HS_D_6,
	output logic [7:0]                       Tx_HS_D_7,
	output logic [NUM_DATA_LANE-1:0]         Tx_HS_enable_D,
    input  logic          axi_clk,
    input  logic          axi_reset_n,
    input  logic   [5:0]  axi_awaddr,
    input  logic          axi_awvalid,
    output logic          axi_awready,
    input  logic   [31:0] axi_wdata,
    input  logic          axi_wvalid,
    output logic          axi_wready,
    output logic          axi_bvalid,
    input  logic          axi_bready,
    input  logic   [5:0]  axi_araddr,
    input  logic          axi_arvalid,
    output logic          axi_arready,
    output logic   [31:0] axi_rdata,
    output logic          axi_rvalid,
    input                 axi_rready,
    input logic           hsync_vc0,
    input logic           hsync_vc1,
    input logic           hsync_vc2,
    input logic           hsync_vc3,
    input logic           vsync_vc0,
    input logic           vsync_vc1,
    input logic           vsync_vc2,
    input logic           vsync_vc3,
    input logic           hsync_vc4,
    input logic           hsync_vc5,
    input logic           hsync_vc6,
    input logic           hsync_vc7,
    input logic           hsync_vc8,
    input logic           hsync_vc9,
    input logic           hsync_vc10,
    input logic           hsync_vc11,
    input logic           hsync_vc12,
    input logic           hsync_vc13,
    input logic           hsync_vc14,
    input logic           hsync_vc15,
    input logic           vsync_vc4,
    input logic           vsync_vc5,
    input logic           vsync_vc6,
    input logic           vsync_vc7,
    input logic           vsync_vc8,
    input logic           vsync_vc9,
    input logic           vsync_vc10,
    input logic           vsync_vc11,
    input logic           vsync_vc12,
    input logic           vsync_vc13,
    input logic           vsync_vc14,
    input logic           vsync_vc15,
    input logic [5:0]     datatype,   
    input logic [63:0]    pixel_data,
    input logic           pixel_data_valid,
    input logic [15:0]    haddr,   
    input logic [15:0]    line_num,
    input logic [15:0]    frame_num,
`ifdef MIPI_CSI2_TX_DEBUG
    input  logic [31:0]   mipi_debug_in,
    output logic [31:0]   mipi_debug_out,
`endif
    output logic          irq
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TOKltIo7Mfu1F3qy7Jd5jJFnHaooxdmYr8ApUO1lRH09S57cVX0+VUFdhEs1WssA
dF+nPiD5BjH6pQwpJRT7MeHYcSyKxD7eoKgTzihp/QpFdBGUZ3WoqYO38JQywc9E
kiF8oB7Ujo8bmr2rKq4PNScIXV1wKBymegt6EShY1Qa8ic270ajpSUfNGnRnMjfK
rfQL/jfhXgFfz1aB4tfQpZdlUBgK2faUXOyp2eWU1chEDiKZDV20qMMmjnhlQflt
/d/nelbiCGsz8Q8oUtPqfb2XMDT2e6gImx0Rk85kX2mG9/DqIsLHhtpNGBXYjW1V
mppdGcTBsXIwuOtapE+cug==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7840 )
`pragma protect data_block
TY8E8kgSj6sbhxpfMW7J7hTXzt6JsnMDQxUfGfC3qP2OCE9MyMzm3reLih06WjCn
wticG7xUtcxUKFzyBTt030GHdHT3+wA80BHvQ+OVHTwTSwylEtQtq7dxPjMGV+v8
tzXhos2cDJrMXkPZKQRM4ziJ4d0NmiXHelcbpVdKPkYeeYaZxA6JysATV5PIwR+1
XoYdgrUwzW5qiCL6qVqN7tCMnXpmVdfadgaNe5SL75CSI9lYg57TM9OO2ZT4nFka
Noq9L6U1Y19kXzmxDiRg5k0y/my7QA6X1BZXh+UjWc8wyrZE75P3QZRzZp2Evvso
95HplDB8Xo+Z0DOOmiQisxtMjGXhFaGo3FiUPXh1WgnIo6vrYp21BXwRKr4fFh/O
LtXlCeM2IntD5MgckM36gYQrnzAWKgbnIsjz7Pm5ET3j+mNENxSRzvYTRgwlstuO
Zl3VamMh02ih8VOc011IxIc+gMtYGM4qdijtLQtTZ8AMjWw3Iao2Xn10DTkaIG7h
CzW68C8jlvO9mMCgMn6BrPZacqtF3VyOZxF1VlYobQimXthbn90EAozyiW2gT9ey
a8Izl8LCHuD2NYCwUkleAxxdwSSt5sBQfshInR5x/cv8IZdD4fkyiPjJC5Wxo3jG
4vm5j/LtgdzuBfk7rjk5APjdEDam3vRwG3K9IYbo7jKFgN8oz8BQiSGm7qCzD0hI
lHW5Zld63D2FK4A8V2XDMGvQohCGJJPw22NXRX2xRENkHAnWJ2CtVu+0mF8oxIve
QsoEnyr0RHu81ukdFKaj1uxImEpmjX//LOkf4tAI2o+3rbT0z4Iv2d1eU/s3Xg44
2fezHrTgkqK/DmW6ZU3KTZ/p/LAwz8/xIrBsyOG5lMwbFCFd47VxCbRfAOvGKjZD
c3dIXPTNuJgOTh/ZbfU0Y1u9IkPL/A0d1mGbOpMppErP3SLdYOubQ6jZ7qBAHLy+
/zNICBNAC4lw+zJ9SI11/NTl8dQGrdu8nhD0PxNhJD++ZmiKdRPeG3Mu3+qXXToL
nIJRFh4B0Mcy1VSIth3lEeEP6jByhSkQ/iXwTe4ENj1sMW5DZg7ik+a8vvB26xXj
ulRxa/DKhToS1/rmWC6MwAObaTOCmEAighyxtMcb7MxrDSls2eqrKAoraF8plgeL
efcI5kF4lhGqBOfLeUtud4t0qV9bYqrQQZf2GvZwERTlim4nFTehoy4xbXZWx36v
8iQ0hJaefgmJMIhD0PDkYwD8Ee5G/fZa+lRYFGQZap/JwzXZaGz52n9sj2zoWx5p
v72tfepzkd/jYfS4tJBQU9LSiRSDr/3A4wQsQmKKV9iya4/ol5tLVA687zJ377m1
P3BR/2bS1NzZmB1lXaoBErKByrBeDsSWIiR06f+03BNA1PcfjxV9KboMTyxBS/zC
w+khwCoQx08KtPK2/9hxayIU0CmLcCy4fzfXrkkG8NI6YsewgUdVR9dNwi+4kNTU
4kzfNhlMH0Pyz+HLKQ3RxWlKEoP7QLyJPbRfvnwLP7X5Jd7CWTk3e7tdFQEX4TQt
sdYbZQUscVLm8AEDEq+ew7ycFuAQNp6Irp1x3rNVJD+47ARvdeFkPpRmZ4hgPpJB
9kdU7CPlW6hhLNXiBEo9wQxFH+nacRQAYMwQhRAM4eTK7dy83IJD+3QYZHmrv9mH
/rB2tHqoAdfJ2TfEOV1R3pYeHKvef+mNH3EDZMU8tBZOwUL66Q27qYBbn8zaQELD
h/88dc+BeNZcoeY122uakwpN5rcECQaz1Q2zRJVJtqgHuKN+w34lNq0gysYLOodK
xVcN3PJwr8xb4aBS7ScBmXSXtSRR1tkHWEbNaSjijaoBvjA5+e5VtNwqOAD94h4s
cmuZ8L56etaaj7GCRDCyeYyAhOpqNGXcQSmQGWJjsMdmxy81kchJYgUHD3i2wgbN
CkvpAsYTLVAGHAreU3y5AQpBL8nYB/quHCEkmCDsiSTNxXAw7aMe3hCQy76096uq
srQG3Bjv+Ln1Xamw5DHF5GXN+CUBFjuVlNOT0WtZ9xWLRvRNXSQVZJO+Sku6lktf
CgV7Uj13y1LTo6m32UPCJd20+Qzf3vYSAKrEI+KYR1EExxHXrQfEwhnHCWK+jYXP
MYXZ0j1K5nkiR80WR5+L/tVydqFbr1bramzAZjeRIIm85wTapT0FJ4gl3/hiEerW
b449xyIGN26ljJSZcCN4cOl7KR4KJW+lgTVLaFloG2VEp7Z3sOKvat5MaVPRyORT
3qRT2XiSQtOIZhuV9tCVipraKCYvdyXKgNCachyHWefzfEr7x/Ed3HaV6/sZmCrI
qmtRCCvQ82DjJ91uCSVIbnTycNx0LqcQcywpEL6i7LEGakPmTtRj1CAP6SrJciL+
QsUyLDWtsdBDpxnmryADvYU39FOH9vRtzWbAcxj0CbasHmkMnr5YTu48FFdLNty2
FnZxc0M8W9lOzlJ7sKaNjItR3Qm/Gucjw2XNeZ70+HDZE3vxPE1HYP8yeuIS0pIK
9EpsO5nVX14pcAjbe0cbXarpbfAI1etDPzAywpt2pDXkLR1vZmQYYPPog/1Dto97
nikpRleL9L4mZ14eYXpwYsAyA6UY7qAstiDmu1uuf6h5RQGPfuZq5WSyF2mksEEA
SajG6EAtduMQzN+S2rWoRBsXNC9Pl5TpVB6KbtQMLZwoIXgisxhzutDjcgmrOWYS
Sr1b+EDVie7O0FDQ6L0M6Wo5faOEIcT/eQDd3jccqZljQ7Ie//Bnz/ZflG9CiAk1
m4SLv2N6nHOvSKeXfPZPxXuxSE4O7G2ssz8PEDHYeXv+PMhs+wCMXfiGc1zoE3rf
dX4JucQfiD8r0/+FAhf7Nuj/HlS/DpSVkicgCmprsFDLsHhRcujZaXW+yRsoJHKR
xvfYGAofmGPrIJcwU1MB7CS6Dq9zlu2FvndJnnuXpEc2dvfY75MyTsrWBNHGrf5Q
cwqouiGbUJyLJeLxNVKFqIUTZAvLF9fl2tFI8o4smFJDfBJWyu8XDK6uWCefvQsO
7HUgc7Ne7G+bkDiJsNieE1RppTCl5koM9324gqXvYD8Q5zm40Mba4zGfjQsumVYk
UeB9kvSKCS4NkHZoitEyi3tFqbX8VKvIjsUmDptVVHOzWrNDrAwRePLSgNMddLu1
37lbClOmX23lNIRO+nEHZoTIECA0vgqF1edsi8bI35zfs5Yfg2XVXFBeZJ0Atqol
eHlZ0MsdZOqbW3MvElzpbON0U0f6U4AJLEm0dOmOv/EOoybd7nvk986Lt8iDQt01
Ys/yUF/wlZf9dS8eyqm/yGmuQC6RcgMgyiJGRdIeW8mLeOvJDtlKG746PL+igmSX
/M1KY48JBVA8lOMD57LlkrZnSseL0i2CHLM9lxVmwtP1i7soX8Ni576Lbvi9KOOm
QjPbPddxgQTgbpmo6xSxCOtsLnNuUIg4WgHTSkWeaPKOxWgZYdSTQJQG3blvU+PD
iGfyU0uK9q8ifTqArTpy9rbSSrBwG+5IxXcRIHp0VgD+hQy4eMaNl5obeOKqstUY
eoTET5SDVIPaQHwFsxlJsYqTeZN8fhrumkM8mXQXBabqNOatugEXovybuQwRh3jA
WPvsHx93xJHTyDI24amnSUW8Xp0oKPnPZLZ/0JzZoRQV4Y9bIz2rMTAObaQGPnE8
CvEyIaMQ243l0kCn0I7sNSyUaJ7dJeHZ9k09iTQ/k4MjAK6KNWKxTvAZNvd2nCCL
Z+2lBMk+6hBACSytVM96tbHVwrvjdjOnCNb/b6lgQGc2Y7pxVfC0tlQJOqqxfZBt
NezNR3cW9Xi94020fHKoS8ybaqMn9Eub3392iUq7YWScAaXByKGRo9/PCbjya9Sf
XHRMGNKg5rbowKE7Mp4iJpjgYn76B/hxjjHahX7MFwJAlEcMemR+Fysvh2VZgUm8
h9B3rr7vScMtFMtp9d6j5f0VDI/texGoqNxDm5YbdxXLEH3dgNIY76WPsKIkGDmX
gJj5Ns+FA19geOnpV4JLgtngXVhSiqilZyn+9EPxY/5SUiWpb41x8VwYGM0AUP0V
fnGReorElnIzEmfPKFaO2B/o1MQ5dBYSbC3djKmB0D5u+K3szFutsnDGStvpYrX5
EPWzhznH/u/3EsgR19diQiVaNwCyMge65DHq2pESOYJcG9c3soLVnlZnijcV2FWh
RVRt+fBvQMVRP1aSoKp+lyqKvveIMB0hzgGNXhoTi5LsGQ96lJPWDDka3yFf7MBw
R3bmIXth//uVZVSAG70ZMcunp+3EUI0B7Oo2R2Pq8jEepXwWnJSjJaJ5kkTmoYy8
nlztQsqjGfDQ1vKkPqQrDvHDoPEqdFUHNhblfyGuNg1QKzFeA23269+CEqxHKRfB
TzOWkmvBd7Vl4Rn/PYBX3dIA7qUFaZzKeOQNegkO6TS9/L2UY//3okftMoHd4j1y
5X2KjUGOYsyyjf7BVtDcqgNpM3jg1p2YCEXthBhBnCxirLmVtUP3cfPRDhF8iJ+k
FZHj/zC3OK1Rz2RHHW+7/hB2oRBEDwX/jBopiwhkgbtn2Bb+nZXlYpo38IqTL1bX
HJcLVw/KPDt7i34a4lUvG+w6kYh+jlwcHflsx3l4X2nuRvVpug851Oxv/P23rUc1
CJqcvLGdQLkjqzIjjWlhuNwcSMqaAbEHlwR9UgRTJzWMjKONOjt/i4BEHO/Hg6M5
i7MMXyQC5F+x/vWFFuKN2z6F+ThDrewHl3Zc9985GhtramSU4m06PxvhxeIegiQw
2TwFMXHvDDRvKW1T5pm02fAC6kS3Dtc6RZ8yfXJOr1nwrh3Ze1CZsi6xNn6/rjtJ
s2GBNH3rkp7yIsBG346iFih9UKaSPz/ZOvM/jLhvjg6erb+Awh10JzYy7IlzSUAP
+jsrxMXOn1MZC1VUwNDC7OWlXXK56xNnhwuanoQ0hxrsARGvW2MWlUy6SHAGWQwr
f0EjOQ96K4Mhz5DUIZsOD8GRztxZqnQOnwlHlZonYQabc72rTX3U1HqBBleVKnFh
Jg7Yk6SI0iXbv2PAqRZuXZzbz7o4TNeHBXNELSjM6DdxvmHHBMeho8QG0mJh6OEq
ydOoQbm1L6SCi/YTgRFo6iqXU3M1CvGTfw2Ia9cJGTqdWTMYToEddfK0PAPSDQ2n
xVl4XmVL7GVNoh3OiiZB02Li28WbgmZ2r3VnZOFFBpLgoFV9AKpt9GdGQQgkZF2+
kkgkxERE0jysZpSmos6kboGdVOEvhGpSv5YtP6Mo0JMQp+UTHfwjhDcjwROEduMz
QEtxeBDrOwuTgE7hWftEuhOXiQAFOdjH4twSsWvlh0OOrclQh26Z+Uv019oW+HsK
dntdRituDYJlxgl5ovdu2VnEtTN3q3F1plvaLk1+UDlu6m/j/yyQ3CpRz+zhQWeN
Quk60szw5ZyKTD6c5ep5nd27kYrXiV/E1Ct5gF2rFlfN84fB8gKIANCdokUPUfzV
jet69uNocPFfkERaJl0X4URMW9dStttSM+UzZYh7VxfFINUNSL98/g/E0h+pLIbA
3hZiBwrPh5wkb0Gv0pB1JJ31tqzrKKkOnGtlGYewYXhUAB4pEfttnTbwcq5FgCAh
ryshU+HYK7fOa4K8dxzzqgIg2Lb7SOh6g+0oFX9H9Hkx2Zl5SKWi8NvYI+uBNYZj
b9thPIq7AcVe5P0fVg+O0dLuh0kAtvbOivQHno0CFv1TfKfQEZbu4nSaK7ne9Cnv
crZPiR96/aJE9bDJHLZF1sqbj9nB8vsJnTYSh6108/ietBbQJGgmYC0RnYt6m23f
ZA7u2Vx2ECJVjQMM3nfZOc4VYKzUr++W3LqTbqheoXxjVcKvkHmStvp2PEv/TjQ8
Xoym36B4/vdf9q2NHlgbR/Kw6mk614k5ClhCS9tmHC0tKFbAfNJUCuRE8o7zZjjP
47POUg8HsUqPUtwGTAyf2QUgjZGG25JyvKwFlUgGf/uljebqDcRKada5LDKI83n3
IA9WcP5/k6AxeqQ32qkXdvg0m4C+LxMiET1lt8ELCMPWfX0n/a/HPh4/JVCPJwCb
W5xOSj7GwQvAULAtrCi174rfzOteE8x5FmDDidgyi3e2uerC4BMnXHcvaCDEtGF7
FQaDMNFLUzgadAv9sFQeHqpz0DrY3q5ALuJntmvpnNduiJi2JQwRlfa+3kNERZtV
hkJo+E38s2dfP2C2qo4KIt6myWt2r7uyF/B3a0/Gu9FgHzCHL55qNf0BooZOOCi6
YUDp6SzcqvtfR9mIHNc49ka3zqUKoUvWgO3+vsKyHMLzeHkXyc08ryAjoxEFSjEy
qG/rZSu3TnudWXLxZAPVBzPyaPDH/boDKreyt+FuOKohTlk9yvJY8hVcY/Fj0jT4
HGJRRKPKYak4CNMfA34tjXLBZnu1t6g5ZdodVq1VMLljtHByQgmZmsf/RbAQe4v2
iWbRV7adQId7jaB4wNX7CmyplH56TrbUXAtkSCJRC02vmD29wHB7dG2oYnDzrOep
/xbBpMRQr4z4fdupp/+kpkTXgmb9O0fTTNSSQHrWCgthIAzyg6gFzvzQJxtjjDjm
ZmTlQhTVGWy6SpiOorPuvhHSBkpURfCpyU1A1RpgKX2bz9CD0FhRMMhs79ss6OX5
xtqXlGiqaXuhH9GipJjDcrIwwzts8vAy0Q4YO4J6UnjhttPBYmENkvCkSSs9ywEz
tT8eD4QWch3CC/kKJ/wGRljhFLrBrW2P37ZhB5f62W48mWK0iBt7TSxZiFNd1Kxt
tN8JQboCKT6zDYsivGYUhtOOxNeDkj9t84d3i9inkkMR+E4Kq7roqiXFCCB+EWLh
uQohP5sUCiDGzqyvjxECWoRmwflfR+YRYLimNm7R452t1Y+tDBaJ6YNrHmYTSiLB
J3lDkLN20Cxxx4xYEb9ywjhMVqNPJ5sH7g8zq0h4xbtR2lTXR0RrWlbD3AZHhPxt
xQ7Dt6w3JSzlniJuIIEhClRyqDSvyROjr3xu/WAahGkFwbrZc3Nx/PZgKx0EdPzw
CfKMemxUk3D/PJyuxLAsNr6DW0wKkU5eq1/tNNKjm602mWpLf1GYxKT645TFDMfw
letokfmXdxXxzm4UqxHI+EyADvic//kPS1HrTQaKHVWRqsOZnM0Ts3buTNb8+PLJ
xdLHA1cBelDpMQgtaiyWs4URXYd9JlP5i40iM5+nAcGmyNJprRtB1SVLVQjQKLKs
4n0uJRAu7AkQstC2B/oi7UZ4anxhw26wUcEIFwvLv88PsVBNcR2s0TAu6xlO1GAj
EA5nyU40/vxY7VGLwiODtxcURaQjvqyQEyir9WTFJ8TAhPk7fa9u8JxohQ4c9F7D
l4SeUldqoPP+wD2giWsT+AWbsC+IV0OC6+nECamJjBxqPb/zAFjvW4WWjxTRnHcL
uMRx4ipIXlerk/kyu0BoDIPuL5IChJCsAu7n6+6CEvDYDUuci9pZCwn7IQlFKMgh
P+Xe5gYmYxyzW5qhFP8QFtpHBVusemlJXOEd5ecs29cJT9b9XpnUZJnrih2WlFDs
6xRDUP5RLsR1AECvjT3hOdUOqtsn1yGWQeryFqPf3SOXcxKdykRyKRHXKrWsq1/a
LuJDcl2YrzCOq8xfQKmTV6F/oqn40fYmJHClJiWNQpV3TeuPu7WAhk1k0jjwbTDJ
/mRLGvAhDX9zm13WP4O1/Pmn0v/upFsqlPJfcJDKXoD9jzsccoJe/d5SvPonJB3O
Xn7AXAWRlOWdfG/5zmn24b/4q3RruYggD5b4ixq4dTopWGLXocvKS7RnInM5FSfU
WNWIrMnIEdULHfPf+OFqSyjotmn8k9onx1jA0eyGEkI+aUFLAEn0dzQRHA+T8jrc
EtozU3BNtMnshdN4SRp+t1G2ztZ8pnHCbSthfYpT+a100i0fHJnKrYEIU1YT6XeX
XI/2Lg5I5dOh63s0xyIktx4DvcUDCL+R3jlkO+l8CmnXemYW2KavPFP0YmsMNHHC
QhdEkvie7a5TPFSWIbyMcS+838kepepbHF27dfaVhspmr1xRQziqIeHXFqdWU/Dq
HqtJ5mukWNdXseaODITnY6bxdYp8gpZVjuvYndiXFzEcwXduMTIjPxhMKdtu2FsJ
Po7oaUWb0Dl+bnUuda966ZA0VheT38FnGUWO9ciwrLswRZdV7lESRElAOrL173Yt
n2LUlOwP1TrLRmXboxQiFsYtU2YKQ/ac8xLI80/ojOVeJQkjeEqalqKAkwziArAG
R8qd0uLF0oauOOr1UtsPQS9wG8S5M47h5twgYjrfDdiw4pO+6v0UvoMCa70Q7GTY
dHzBoCZS5FH/bB/nbGuoxjX6XU6Ntb9B5G/8Bal+5ZTbmMFToD6Rg26oYMKGiNoy
RaKWPahtsvV9qYt4Lgxi3ueG2yGxc8i2AqjOYt+0B3whzh/XNv7WCDvIoz/0W4rL
hzTwX5yd/5bQNPznq0Vj//d1LA6+zIKqCfkIViMO5GjcCttJR1+G5c0oWjuL/wGh
Rgsw9MInLALQdsA/M8kPeyKHy5JbmfbcdGCfdNF9cAdc6oCCjIWFF3vakKvdX5E+
4aEuCEIriWQ0cYNXmTrvSQ7O5OYNNicSlQUvGjbtDzp+hucxSUE0pdIuugK7nc1k
CAOWErEAabIJZR+VM3aVQ8QIe6oLDhjY7JbhHcw8c+0cJd3IhcuaC1lGo9TjMGcJ
9faPhysyVLWEPltVrm5diKyETezVaDVf7L+mODdFwqN5IXmoK8lS6e7JZO31sIXC
QD2EDUTuBJwF5MiEtYaxSY/aI2UqSgrYccPtY3b3JUTXCoSZUSTiZ+fIfhKWX1zL
kcy6mRaLUzSXzPnej/s/MG21FcgSrqOXynd+4EaeUSrXx+lyXW7EZXSX/rYIvMmW
280NDTj0X/5ou4QrAzMDgNGMiOigafnETICLErUPjWzunWLgSrbCoZBCn0DZm7Al
bnIBdUOZqc9suQHtjlpwCoBz0VEjpfTYFANh4eBJQduhYcioneQe/+lcxatfX2CP
lH2EqFUQitfD3ne3FQmkPNCPVfS+8dJ601uBqtnsGkoSlV48JmoAXpkhsy43l3n9
xLCUBZAE/ZFHFbTgBWUxImSw5NKi01LORSI6j51afwsTV0/90DzO9EACgnYNl3+e
wVDKoXsGvSFFtthbRtsrT+moI11eYkiQYCz52gweUFV5De5gAyd1NsrTPSzJSoYf
okTQyZfBWNI88fBEzMVMWhbIDfGq2Ut2lyQc1Sh4LqZtk2qKX5UZkbpAc+pJCS+w
nmhOc2lMDg2o3DdkmaFg/Q+Ovd4B5ZMX/xOQRLKpL1n5xbFYJeMCvwQYQChwl1/I
CUGXyurSmxlYrEz4FzBGBg+61hDFsNunJCNA4jMrsu6fGPIE7CGZ1J8dugzKWro6
TnMjZcTlasBnYWwf9/kjFYLS9iG5fmCFRU6KUbOdvEz3Fx/yR1twW4UNNUcAXjEp
85s8/4nmWJRVQf37Zqfw1c6vBOvhs1i0tUefCQqRslh2hD0zwX0r3bvmvdotXxy5
H7nMUlFqiwrVic1YcmC0cfwSWs4ZdqAI5tOAYk1OgY41txVToj0t/bFYYuZr4nPL
lUhafT8xG5NMXTxWgAf7l0dKjeE1bMUJ7o7di7Wovmn5Q+4ijkTv6k+bIpKZT9rt
TDO4+nCDBg92DGYr2EnNzsOCa/4WTOz46njdo+zj2hYROyc1vKiLNntMz06fa6za
PLhVsPKvJMO1THHjOEPcq5wPZYVaCPLiTU3aSUrHaDWQ0/l7oE1MLwC05hmiqBDO
PrSyaj8Pb8xpJ848M0DppKANknMhZEWujmZ2kE610KNcujY4SV70ohioykH6i6+P
wT8HAUVxye0nmAG2LWGOmkhWym4sNshxT3eYoYF7m+pFhu0vgG87MtJxIKQiHy4I
qd/SeILWZog0jFCS7WbxRKy2pIpkJUd2vc6p/h6feRaduwhCXDeMKznzymCu2ZUK
/2+E4oufFy3UQvByhufR5A85puW/m4rGSBHTt2b5wCHnOKhTiz+VL8TwAQN7vWm9
91RfiUhzFY9zLC1/Dx+YJPFDOl5+YgrLqK4LZacH8ggAcDM5nc6wab5sk7tagTnO
Oe7+DWohxoxZuEOnwc7GYncYo/sZfZc2CvdpoNND3dqP2HV251VZMuZ4I+98boP/
9cPDqbL1k9kDoKXME0hfUawZOmqmCeCkwbrrPSoyGm7lKUGK1dHaOi+steqfAU55
MG1uNlWAGL/1H/N+XnVW0UJ0qsv2TuP6LcMjUc6nxpyiSDVhBU/qyO1U/3Fp1vAa
lWpLvOwgT82lwzzwIY12A3XkmTmPbybv8hRUsdIgTzRrsv1kEeIrpteYJVNagUeZ
S3OTzoFaNEYDH+q/zkijHQSxJriKhFcm02HJaUIWhxNmWuwqCdo54B17JwwjNYa9
e48fvKZwSbP6/3r+TAnBDimQ3n6p2RUmjeEpZjn7JogC6d+VRxD1xFjA0pZNmZWx
wugnXNJbm7/8rrqOaJtEJg==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lu2WC7gBEiAtWDB9o6DYPXg8NpFZxld77WXd3s/S33EIIEk2Vbfees0rGfbkM4cZ
bBVTPsZqpheo/5vXRkg6Ue8efxBDIX+KIkkinKHFAFuOhzypDxlqVtv7QH5vPsbb
zBC1Zdt9LKk/U1ItTIAN+bZtLcAGznMJ+yvB2b9mZ5cKH5b8uzYMQ827azIcHFf4
v53FNd8SzCfTLc/a+YSC2NaKVPluOeEVgqsikk66BHswAsu/DrLNNdmJRq0m38Tt
7rpyGIGpZLUZzG98Vjunfleb3kq4m+FgTIDlU+ida9JvyuzaYAUKt4GkJJByaTav
gwMKL/3shNDfOnG9KqrTSw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6336 )
`pragma protect data_block
BIoJ7jemCfHYR/fPV1se3wg9VmWCcD5xxqbr3ta6bLTjisYfhLNrmvCRuAirA3xn
M4828+o/+mA9UPPaXL4+0wyelH8dwY9bOFtLK718WiATUQCuBdfjPR1Z3GAzuc6+
TAqZItY+d0US8GqQHD3du8PryaifeeqOX11TdsXifX9Ua6IpfYexwfabbhhH3rpR
iodF7HHUY/dE+UrN2jS4BwgDc2QBHBfhS6Ktxb60LIo9kv6y0pj9De19Yh7j9ase
W7bCEmnVEceZlCG7dDRW41QU8P9B3QVx+LdlVwkPjA0sbIGKAw42mH2S2CQMalgI
DQ3q3WrS6OsUrZY46aUiv54TIhYDXu1zz5LBR1X6PoTepuhwa/NhBGIbDEx8TAiB
77npkMx4XbQoHGsXcrt6g74NaPh2nK1AL6905wWBinwK43ptCeVZhshM6vjHm0Dz
az4VS45RYH0lxGymtTe4Gy9XZ0sNSUr13EdLAq8/IVs5zwOiKUWW9EwiN62oHMWx
TUzHye8s2hlObfWrjIW8g1UatZ5uTQdAXLN3/RzTsF5Obfc1TbZCqX9cFzHddJwF
nqJ3n1LkKa5ZAtbtkxHOI1dxIDT8AkimGHlDluB6JW5jyYFe8QNLbr4Oj6ss6iOB
tID3mWv4eKudyXo0BEvTWKAkZ7Gba9s6BhjPEGq8g5EMx3t3Dr/KBw8KSh/DKDJl
ZiqNuBvvC4bhDIWkPp8zLiBLj5C969vClVmm6hLm9kPfnP1Y4ocy63+6Tf3M+hhI
5bPKVW7fnj+3UbSR8LJ3pXEMI1vvoPruOB/ZwxVYL2jqJQ3ypUCcW1aiGHfhPwlk
FheIvD5guaWNy6lzVay+1KHslHt6ddBE0CDySXLVOFcDIxEdEQfss/XXqtQ1STQi
MT4xTvVp/HRjeICG7MC6we69zntG14se8R5nUQaoi9hfRFoUVx9+qbjvjzP/ijGe
9l4khiVi0e2YLz245+E+X1Mjipz/Vz63Gi02l3OWhb5BUPm1nhj0otXCRgXKonCk
r2HaSB+rb5wsUWXzkYJu9fiGHeyOPMr9qenYLR2OkY5sBIA00G41dyBp+sAAZfnN
6tnRKc277F4aOrZXC+JtwFeDtmxnhFgowpxBnFn9voZjNp3JRyXIaXpwPtcxBisD
7iYwkJa/6Yx1zO5Q9ddHJxGVM9zPDeHUvzpSqjeYDH21z/O3lXetNPONzxhy3+mw
y8SEIixue2B8zYm70zpOLsOGgj+nP13K/XGwqtZTc22vbiI+w1tSNwuNY9ysQdg1
7vfJLgIka6p44iVe9aHzNhAYQqLTHmR67x1bZ36+iriUWSy54dcVwyc6yr00PVBu
ys+x2KGQdOZHw/ZJoZHNYoSC3f4yFpNLYs4rrpdmL6kf1UDkUvE2p1tilqPQNq1O
gAYUKAGlob2hYfAbqYhpDU/wx0UpIvR+qcWcwqvTfrBl7TVK8zWWrpDLk04K5u4Q
BHtNAEXypbMIYnseJBKcCgKAT5+jOSqiuchQVYPooSDE8popWI8uQWP7PoNbX6xf
/4BGra99OvYECGBeOD6kuiQ+718pl8vvkdKuECYUzSTdFJlZT1M/UjXq/9wuNAuK
CM4Zm6vqPJxPKlEPARkGaBSiVIm8OCWEZJy7KOygxoVW9q7wSv1O5JDeRLH2818S
OsfOAZqirLCm2yP1GJydHIL6w4XCTHJ0+OX5+TTHe+/WIm2SLQQd5c8Byp5WqEPE
l/q2hFhi+ItiVaRFm5xkV0mwUqj6DuDRuFt2TuiAnLpzmjNZ3h2jIgQD40PdMMp6
C4eIarpeW87ppWz3I2wGs7HcWytqqfTuK8K2f74XnZSHHWkcupX3I2MgZN4SURzS
HGwfLgWJ5aoIEecAwd0MxbN+el1Ynvopwthwf2xquRazTfkEZPo8VllnVG6M7Xki
UjxRVz41A2WCFRjVWoWt+6VBu6csujCcWeH7DWPqDlymzx9/1mJKvnBdbpTfA37m
7R0PG9Wz982R/C/nv3EfSP1TZC/A5jNZjzTLYu5ZMhL/oRivM0VlIVOKCwsb20bZ
xUwsQW8VTXqC+00+Uh6997rVtdeshPhD3pdnILh6SwLIJe21ZKkQl+UoywUlGRu6
QmZznQ/TbN5uJyN16ZmQTwYyt9wwT0hL/wZxg2RBHdwO/Wpzx/HE/RRRbM15f8qV
mOBwzEcx+JR6oDZTJPAPYjqcAG2Aj/UUwGUcWkZBpNr8uTNXi/0hWD5BFTdS7H1h
f1FdfcYnb6ol2j/ktvDzBPP9f8mYKS4KIMlGj3+hgdG/L9C/iXZl2ovf6ooiqKDR
c/demICX+HoeEm/as8wRMR2MV5ZBMtuPdELAKG/Vz621JsYMijgZRt2c+0hVq6Pi
RP4f+797jH5kTaK8GYOaihfw/P/cfOHVMmNrct2su+OTzi+1EIPk/uf8ZdtXnnHw
WfvEcWhxrBUXd4n2YZy54CbRyseg43SdEy/9XSkqbsOiWL4Qo4wLrQzZwvcBlEbS
7rSN497H+Vob+r/85MTVEPhd4MujQxVsbHqgduglhCoxvh9nvGYZGtekNdmuQJac
hAbsQOjb4BldSy/LU4wAEpg4bUlTQ8IsMcJdhA6bKTdB/np4kFyyttey6YejyqNP
+Dzmv4rTJ2kynJkCoS/2CBAJmOZVd2f69Xl6FaG4tAPBuayxD7IsAWpj2b5WmUA9
wYgzZeC+Sy9XQTzILVlGHn+rucUBrSt+86yZqA0ec9hyt2c8VbOYujhMRsFZFck+
NFSalRscgpRDqY67Xm3abZo1dnLsfGpH5n0MdhJ2COkiISp1bDucmYxrFSCB4PKl
ezKtjJffOR4nraY3Ssu5pLSuTHJHUXVZXtrCemEcgfHkMRWCwJlprmgCrdNLeVP7
l7ZpqgeWDLvzJWP8Wc5yhGbxFcJJZ77JXLsj67DXiBczYPme/ysgMyksT6KxgEDd
IyM2mmDF4wvGGyraJnFm6p4dHzJuca2gE5+Ib34zcnRdHKgy7R74RCmTstFRqpj3
lJOzuxAKKawh3yEPxycNEXEq4qM6MU9z5WIEEUuEQ3dtfX6mrxG2Flvu2mjhJsY4
yFpz1FL0Pc85KKv4SDG49o3bW9eki6jWnW+wnZTVgBYpGFaS0uo7pkjKA+e4uln5
SpTUn2pD6lWqrQ1c/VPK0KytURJQr9pgh3pMrDID1fdLNrH95bDWALu3cxUXd7KS
x6HR29q/iQuuoYgYZetJEwJKhrnNbQBwSyBGCRFqqy/2Wuid2/Du5EXwOeP8271N
Pr1IOeHF8HVpQyebJLo1gmkQXzbtpQWTNzrjjYRtSiVVsBsK/O4e6pXKtSI1Kbtz
DiTrTJ1W/c6AHWHJSjmvOE+qt2DwozxU0fcWHj9Vv81HtuAmmGHr+kNNNhByz9yh
Nk0ziSN8i0mZz0+9mzba6BPQrQkIqERYsoIVBCx2CeXnRns64EplSVbM4Xj3IF2F
FuQkiT8DZt8S4/GHZzPSvmT/+oicIWtzFivcg8ZHukv0DdyC8nsTGz1bRzOu04E8
eW3qi3q0ItI77aTIWyHenvwAxuZm8VZGxk3XKAO2SJKRGgqd6yBHx6IQWvtfu2k1
IYJN70X/3BTsTIC2wL5C+ZOFlZS4V5D3PfEiKz+WYgZDS6tYcD7QCtLZn0y+LblC
rl9Bfa9Wi87365GtmNOQTpUk0VFm0jzEef/XjF//96hpLfog3MNWuhy6P2tRibte
Wy7qHLQC7Qqpgiu7RlRhfSylpl4DRCudgXWsX3mo+BEMNQfwrotgNPl7oyVCYYaz
pD3XjF55aGfHpfuwVjBwHZGs8gacOYtjRxpngmkjcMknCGnRgEsZzV0LkPiR1FwJ
yYZx+NDZUo3F9g0xRmikLHoBDQ5RV4Pl3f5yZkwlRMC3qTfm+JgcoNXggPefi4UQ
OCEvKNQgH7f3ekzxj83wwt5GrRoLFBdoZnyLwexqWAkcvVUG0+H3IkgrFF6uODEJ
BP0f/Z+zIE5MOydcbT28AnK5gDJAkmsUg006Ud3YC5F/oftV6tAF8QpTKmVkgTfM
0rdMZfFmAIGRLYCXsNHcQOPqTKkWBfrJRhaWB8QPBmqpGB4gH89hJTfBNrLz/Nzi
kyj2Y7KPaKAaQ6z50Lh1foOQgHrIP401y7GHvh+r9UDrgk+NhxvmYyeCc9CcaHns
PskPdYltmaPlwCLP0dck9IZa0uGN04dssCijMJkKIoOSPwx/vd16YxdMbrX+YB8E
J6YyMNZoggClWouHUCjwlZ7vn7EuB7PMLaurmZefchfh3EjoxE20cJ7I+mcj0ogP
HPf7G9D3WofSyx684G4VOJsCMdtxV6TLJ2eoLbJtUCRRsvFSYRpWIrccKMToHRqL
Bv0AY7LOhriMg1z4pQekGoY62tNvihsK6yG0cCnB8zNeZKKNgiQoH/DkpilEOiEl
tQgWC0ECQNxA3YmErkrkvNJl/IF+e6lFm0KpFZ/wWJDW4Knhk1+hOF7/gFCicRSp
Y2toA0fGq61PzVBUT65D3M5JsvVXvzigaS+8J1fQcTBxq1c8WQJI4B1+1kiQzS7V
GTARL/4bOPi6ulqeDfVd4epmCNF+10oGcDSozKZTX4v4O3V6iGzwzEn9MnCXXe87
74k1WkjjapQUmkMIdm/IR4gG9ca8o7TaDN/Spsx+wPmHGg82A4QXPwnFWDE+cOoQ
3ylgbHnDZVBspaHSLRr5aK9QF9L0PSgoo5+gkCZyqOvaxBd1hUXLXdAXNPqUCXbe
IzGgsTpWY8wNM+LPVc/nPLggOhBplPzeodqF9rpXieO2Rj2PWfyLVgDVN8u3Utb0
PeEBQWnqXNZrvnjcEQkuR72e5O38w81VtsFl8HNGRQBN/kBaB0kZVZcXvwyoYspf
ed4VU3RthUAsF+SPVSAKx2zZ/hDTG8Bd9LO8nGjU5SOzG1uNrhLL3eJ8waNZOz6L
uBNB+3XlJIfZRJyBT89Um0VhruTKkacp2kmZs/NYVQi7gvOwkpfgmEUGWiMr57Jf
hv2kN8iAxuU++8vsSJepBCnT+J14ctUKj9KVgHng0Aw2azTt6Y3yu6Em9Zaf5E+v
YlXUOfGOMeG2DjgZT5IDjdxRAMNGZgFztq3OlsUaRrBBYCdDjUmuYh63tZWcJGHh
dsiGhwGec0mEZRz5/+RoV54h0gzq4jP0yZ7oaw7EdjyeG/Xlcd7yIaShphQjnXQP
HqXtzUfcax/z9nsY4eKGVkZWk/T7SunQ4Wq3B8Bb5cG0Wt0+dXdlI5ov76Dbpict
sjUripS+djls6y4pKhy+z6LGCl+5TtGqqZP9b3e/Z9Mnj4PaoxwnRotWt8VEiWWi
0lCqneebyGaSZO9a2wRI24LMDX+HYElSKN158TB5173VJDXa+EOEsJkmrJcyb2Xk
7cFoR75ib/kwrbMuznC4th5QAkuGzvH29ddycCTCe1aIuPjCdSMqfWmEGAyfg/Dy
T3NgKEc0W2VGhcJzcaO4sz58OGc0P1qq2KanV9PnJwZF9PLpwbBbfPHpS5dVSryV
35lREeAS1HFGZnGo4THo3QyD5CqTThoU+4UHzmUuSe5Tnhs1aZlRd8piLXolJwcx
oqnSyjq/d3o3927COI5lpg43p1gkdrBm+F0xxV3raXSTu/gkpyC0XhiAAiG9rSo2
l7EfcZoVmSxeadKmvWXxoOy8Uegprw6RRo/060jDCiICM39iGO5/g3eCyu7l9nSI
+Ggjs/m0PvKHSdn2Wb8BPd69yTsPOG1pQLuVtmvYnyn3aFcyJoPnL2SPdo7ROf09
cxylZwIz61bmRdXYceW9u7tUREKtbAygdP5eROhW+yf/uSOC8BRB+aUvseBP2f4l
gwIVy1IIHy+8BA4s6tE4B1mjZ1tXxZQFeNhYUS6JfJoZZ7aDvQfDuWEg1V5B9myS
XaWHeTjf/lIka23hEt7GQSI6twC554GG1gCO2Wq38uq+wnX2RPeEJhIzU0T7jIsm
ZccDBDalCmnzj6xLuhf/EJ58mAsnDOna8jll3clxW9slj1GS1makIIGUnxnHFQUO
65vJuS12l0gPw4BZ19m/R72g+NkCjmSmMC/3QB7FhG5Bivpw2UKasuEleKz1cp+q
JyC7orF0KLWDVdalm+XhaDrujOpCkCtUcPtYOoQ1472qbXz4nZgXrK7V1pUnxnoH
eHzo3ODD8nKbklOkEwVrY/pG+YJlLsfHyF9RRBG2N1lCIiZbt9jD5l3g/QhIWDF9
GA6YhSbmBJuBlFRk0Gqd+SFp4NZXbdiPwRxNLjg9GEIe2PcVpq9enZJCuIpAsatc
ncuDO0cqL3fxuyb243frdDKCiFCgN38NxY8NE2Xs5vVi31GnARYEhVoFomV5GgCZ
GkCJaDSgmRzElu7l2eiLom1ZDopRjytKIaMw5v2ZpN4VQUTh2VQ38Tw7JsQPbsvy
Tt7xnEaTq/fXCTiphf8WZcvZITlswZXIYwxna1B53xQcDr+J2mTRm39f2wn7bZ6J
tvKrx1ZnGvXwUx0wkRkIt5rtmbVBOjVUIqjkesYg9A0ZTWVhBgMYjEDxszmSIJbF
reFheyp9F3v16OVoTnIWjWL/jWvnKdTwQYi4AdCWgvKbjBqQl9+tvg7JxnC5ILcM
PSgcQN/u5+GwJGoNUAyOijg7guq3myoV3GY+R7w858RIaoVskTvIiUsa10/UCYg7
V27vKvoHYgJXYPjnMzaF8VNrWRpIPe5Q3elqmqGi9yKF6OuUhetHdAxBhsWjjatp
06Dv4YQnVErFNI1X1V+u6KewVgXHzrOua1EHsA0gN+k/brjPyMKB85/DlndrDumt
nb7ikjJ11mi1GWw7Jp7bKlRuIxijJ2cOOLZ9tvD0tdOCMvqCda6Iim4+21IJscKu
hGMf4gi9qqt8ObOzhh2bT3+jDh87meYZ0mYNhMlEZl5vociFUHqCL4WSNTf3In/1
a2kvpcTogSyYKhRGgHTJICnKlkpaTpRw41B49VaxYaRO/R6vcpdo0n+owt+oyJNG
bJnQx3dteDtBLAtnvNXV1BhyDrqNPjWgo2Pam9Sv1bug/W38RzmMJH9LaNTc7j5b
fid4bx/bV9gb1BWdCFroXNRA+SeMjd3znJh1ylGKRdVeu9YAXGn+7f5mY8qNqam6
nN6tJijPMZlKUHMWONKTQFugTZYlHL6S+kUslrxl+UzeMzegQUYy6AnmH6+hNBNJ
hT8WFo9t5RkGTSQRH13eRnYAPhbeRYs+NiDtpLSvcoSaCtJdIaNe97BXvLPZDJmJ
XIDvr7jdbQvbuinTQMg76tuCri1//0gW7KqeJZ0wlS0W4HWprIDiXgNkByvboLGi
lNUxOKeUM6GUsAesfP8AWFuT8n42p2rMNKG9lc94vhITNJy0m0lSr/XPBERB6mZG
c4vy9dp8ItV+9OfWBdbM78ehJ/z+RvBuVa0nKjdmbSzu1RijD7ZCqMm+MmtYI6Qn
MXl6cOl8feI4SM08hhu2OB/uMg9tnZ0UJB4N9zc0Kr+EYmDLPszJRZfYeI+8Hu+x
jfOgksiHsQYbmzCGgRh30RsP9Qvy/rsIXMTTSr91I6ZRKIjKxRy35ho2qtid9+iC
Vo/VesmbO/kCs8C3fLGIaUowjyjNRR6E65BiGVBcG4v469iw8tv+/AkpC0gnVU0d
CCg5xNly3RMMWoiMmbZXJDKQ1qmFbQKmw9A0tyzblD3zJbOZcBTOGFB5xG6WHnz7
mC5tRAeijTZgC5IAbR7jRZwbrlJDfKLYGpXL1gEaDoChMHSt2jq2boUrLO5xpt25
aq4aQWmHKjVu4jLUc73zGQsDYniXXyeUas0g5+EYWOTuBBSZb2Z5agYlvA2nsHn+
WUAArnAMKiqNzag2gt8+6xdmxHL6BotqA9auciHCB+C7BT1ORMoLxIpbuXgRUzs+
fd6b7ljJVhMGqM74wgYVpsxc+x/AEFD/A1voNNVKoRMXBKqQTdUzr6d5cCoxqK1r
Hy2g9MTYi2/0W9d7ZPbVYVj0Z2XzhQ8u84a7kFiwKMhJfJLm7uJtfypg8rFUorNi
GYjYeANxAddRAm2tXLBko2XD0U5awPFYx9+b5TZSKVHXd79PV+/14EioyDSaaF7t
+yoQPkZ3w/dG/hZT5jdYSasY/LVgUxwt67JZnenUT3MiE4djHyCh7UuzeMgB2kHx
hlNpP4eRlg0C/gOSt74pMuZ6Bq+6injjFFSj7RGVlLZEIgLxe/tWlSsVCsfXgYYV
PPPl2QaREfVweXp1Bwij/KX/Bg6FCZuG5F7AvhtIXUJXZry5Oer3NzwfUB/37+Su
n7llG4ndPlLXuBXa3Htxr4J0e+uhl2whUbLvhWsoadQ7dbLtnnAunVAP2/lxxjwi
p5EE5+PjBHQaM/z9v5QRpjW71n1mIun+h7dQNGrmMgIUCIfEzY7CngfcftONQke2
7svddvnj5VA4g7p/JA0NjIzppILeETTNaWdKRbuaR/hICSbovp/eqQ0wnirIxmFl
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LprGxna0tDMC5Fr8eBTJf6Y6HVz60C6f7iwh4HbqrjlElOyxXmEpGEjvOnSSxlZi
60QQ5rb5Uvez2fCMeOggJCDgy6Txof/rCfX1CzMRw5DR2QXlgXGtkTyj6fLZkS/y
ByNPcFdXmFmaI99T6MlRBm2DFdoYeWKhklXuoU58JFMNIn2hUGL02sTOuia/T6fN
V0OcB7Hs3xFKYao6xk3zCroWDg0ommBAjzjfOn6tO0/EOMpfQpKEHbf3mmlBe18o
GCTLr8EwE/vKymlOWxWijyfgzmpYCusxZDDOWrShynj78Ul+e+W8sDb+vKtAE/jm
E6odXB7tyyA3+5RGn3akyw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 832 )
`pragma protect data_block
PWpgPjJyBqu8h3da3CgqYlRceJ7ZFlgWd4Zh15k283aiCjFoa/DZR/sEuaGi3kum
bU6tlo4KITiGEywZOPenJo92ji9b2raWzhWFmUE3XNzdBO0C7V3z9rheARbf/BJ7
uPRvX9uCcJ+fq8iFLbAWDBdZM/7nmS4cDldjcY+STlNsfJ3uknCdaWwAt5q3R5Qc
ab2q/FMVoB5J+GU5KPZms9QrbUWde9PUOKp3H3jMQ35rtLTy5YNWvdicGWeI912t
XBMeOzE9AOMNlVirIHmcLbdQsowXnMsgosMHBb3jyJ7WUUWwlXioZVDM8WGMTTaq
lkR2pBu6NOFwEkcFqueqRtvjv26maB9tQk4NG7pecrabjFTCySPwGskxBGNBF7um
+oKrCUzxQBaQ06S6JZ71Sr5k5QwudyrPg+yrPMiFvBldG58qFzO9UIdPvY59rbzy
Q+s9Oy9bwx43ZsV7GxF74Qt493otHPKQILDs1uTI9DbQbnPJUxEstf5tIX44mQVx
g8U8LRPobZJ1IFmZSto0hUOFv64zG1gU4qRetpGjW/sOFzQm0FumIVLN/5bVb/XI
qqZbU38Q+KXXSRDsJA2G+7cebKJ68nKZbXWmr9O5AME1d9MyU0Td9taZvRy0espP
HKJdU8oiu38+r1IsyG5RHXzKMUuM80Ke5ShEdgnXKWvVDKuyzhXTWlg8Fm0PI1h4
Du1vTNuF29pNWrKLnamzwP0s0U6XUG3d/syj8rXb1ECZ4PtF1C9hWt6SpouDrRyn
bISkX0SmYZ+oEjbj7b19AmA1tuYcCrq3kHyAgmCgN4RpAaRbqtKjXu7NlKyRDFO1
OtxLAaYhgFI7nCSKeo/kufLKzvHWuC6DWXTbIKytaacD4BkuKH5XaZ4ShRZr6OSS
rcTHcFWJFjkBZ5Qi7RPQT7nsbKn/3CHRZjbWlsVUzakyURSGSxLQlB/SSEXuHvKk
32j+mfL9tEvE//E1O8oDRDAL+nQpsL0oLbHSnsQ4Cc5tqW0y/t43xquNcr6bk9Ca
6DzVwOX6foZbTn+92VpEyn5rihtLSgo7CcYXyKRM/GSJ0tc1yj04gPKWlG/hf+VU
PbQjaNEOtaH8D0o2lih4Bg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ejmnCX1RjQ6z6YAHLy7t/FREgR+QFCWub2Vb5ZYDCRo1arnvjmUaXqNjQbkPmK45
zJ0df6Wp3jTbNE0SUa3w+SA1ja+iBJBOr/hzkj0ujq+dj88GBKZkGjU8IdGel+FV
rR6+9R5hcg7zfvTmL/BOrGz7o7UB2MAFkDD2DrsHHFqMSstNjt+GM9SC576RRgOH
lVS0sc5JcC7pCS/+VJsLFhGP/GmjwHrcklva5Nb/VFF+3hJ454zC85fbJB/Ziyj1
9Jdq/qCUy/cWrKbE2Cy4cRxFQoVu2EtzE+GcY2Y6vPktWcCZgsCF0++KhX/HkhQm
bCLxTSXpzNhGLFyzB3t9UQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14000 )
`pragma protect data_block
atXdgl2hG5B1IY95oMI+MTVJtf8zp7ZCHSY0sj8YKdiVZ+cUxcrnqVYQLkSgYT/G
ZAMvqDLj7AbRAx3oawGa7YWEG6X0UWdV/hjVTG3Hi68fuYVrRPBZlt3BqzDU8ntF
pJHiLQOUMnGRCOMYmEY8cgF1VtihMHdfNNqdG0NPam6bmNuqi5CsddP2JBirjAxI
vL8qwvFTnuV+VAK7T2oC+0kLCjk1PNEVAlRyII5b0Q5ebtpGFoPId/7VsVQuU/nE
bENyQN2QWprh7DmVCd9ll1gMwqhyQLBuPYiNaovwHq0PvLDsxVDX9mnnBr5WDOuD
jc/SyNr9wekncA56F/w7KpDal3HjZ/BBT0L+y1Yl65AKVK9XvgyREimN2daF86G+
9FvD/8vuqD6jtMuV7zS3H0MEpN5ZAJeOKDbOqlEdKuuOoqWWNrKorVWZ/7h7f9sW
TQoc2NOJwdVMTG5nOii3A1Wqz36bJAoLw6aCkyam9zpOTyWQWbhjloFPiLUD396f
GsTu8L+tTlk2CFw4/o2JWrNzuqOSmvhUGPu8lI/urMz/ksQKdez8A7ZOmvuJYaTY
4mwseQuer5AoyKSH3lpu4R150AN0Kuz4hl4bYKvYecBjmXS/CqqDO0X0Sv586EPB
vn/3CQfPsxD5Fn0U0F1c/IP7jGEK3ejvCkKxHf6PD8iGMxsuBxxiWacty3hefdUj
blTGz2+1fwt2aGz65O/ZVnluzdr6w3E7J+iytsyJBxv+ZZBqJJtDSKsz+XW4fX7e
AU8HEcjmwF5bH6sLOXUx3YX0ME2kiUZ8dS4X0Yn1LpRZWOl8uZ8wDAcT9jrHL0nR
v2RQAjmqlFHorDM4+ph8VCUcpnzX1pUQ/f3s42P3lcmnEuRaulDm4Hjyd6S0yB40
c0ewAFTlmCBE0ibV4cfNYgN43Tan7WbKawGSbszVzHBjD0c+UpnRnQCQ30iilIWL
vBMzPfmTtPqCFJAOSkYLnzWAmLiGI7bKaaBQysfg76cvs2fslSa3CQikhbN2q5Xp
901xYBDSOaDLhqBV+8CgKEtCiMSIZd54Y9kZXzLnJxymYdRSJ5+NX+B1C1Y0HnPf
p/kmeNzxfQ7ERJ1ig+yjqx3iDIu3QGzqFNEn9u+DfqwClo5eH5JLTiP8CFOxlu1Q
Seyf641ZQHNur++BXBHVOMOM1moCY9KytulzgFFxtTReke/skSo5aSOIa9NDf5Cg
UgCboWr74Rt0dZ8A+mF/LCBWwqhbTnX1Gr9Ca5StlRZ17/KO3AOZQYHTCXJik9Ba
EcxBgT8IH0tMbBOFX3XhQVmY7dg5hP72Q3EGZo6319H8QcTJzuvdfpOpDN/tu08+
8yn80SUSRX6TdC9+bMgz8D72lvu7S+Ur1vItIHV5+1id+dfsFs7GvEJD8bH5Nv8A
gIA9WznfdR/JMOILc7dkZul8Y8Hxo9SRa3dwriGsJNyWCHG7lqopPN4mKCPvbyIl
164egc1ZeHo0vtNtKVns3J2MoAMvqifA61f0039xh1+2JQPwIyYyfCrXvHL0vRHi
+sq0C6o568+Box3cUSIg2pQknOPwzTPNxUTevq3nL73jLwnYtuhNJhGpFQPq2lkh
/rFfxztoGOw1An5EkMJnmM0MSnAB4abgRvse0Fq22APYi3/R05VY2muBj3LqRI0f
bls5OsfaJH2gOK1+46eIPRYkmbzM4qWEQ2KoqIcoHf+IB+L+3TpCImzZ7mle0vbA
3gCSuM91PUidjRz8sF2epirsYPpzCfbhWHqbZKnwUT+HwjqpxypAWtbNnUkjpKnz
srOC3llF6wFiHJ33nqw/HoqwjgVeuOqC1GhqraJulwp1jggRtkRyw11uw6Ha5m4g
RJPXKAVkHDrd+oFeQmKWCgcQq+ojAcg62ZrTGDaYLIFWl5Met+N+REa4SImuRWHj
8QZr1PoykmghkEkrxTbnzlKOnZQJ4Z5vIR2qLQ37OGfnpj9+MghV10XifWgAC0PJ
ZyriTUutPu6qVtSMwl5UYoxngbOnePsjP7D8gR867yaBBkibzDnvLP/91XAef4P0
B6u4qa0NBFzawEPNMg/dEeSATEKMXtWNdrFe3OqaHc7dowwYC7K+iXnzGiTzxgF5
vrvCtroInJjcV9DYh8u0TyaHEu1j0hSb6QmUwxkOoJ1qh7uGSuzZByBEemEto/kp
DRY9MmoMpVRPgBYp0lpfZLXYr5qDE4S05iJlbbzLIqBAkqbPftlf0/h+OJErCfC/
EZSw73hXtVeYAZliNq6UqB4g1A1S9TRq0wM1tJZKGjtjsWViOzZDH5Wt52K38Qhb
F7+HvHDxuWp4K2iDZxYqozniizV+15BmBSzlSVUkhEgJcXOCJerBVjKVIW+JentS
Uv71WHLGpgiOyv40N80Y547W6iJ56VmCengBXP3DBnx9Ry+OznOsQ22ojOmajkrc
TO/OILosoIWeAyhYtg9vDo4RTBVQXbBhh14D71ZyLdYCkd0xxzGRBLVcb7LK3ENS
vpHu1oWu2/05XRYLikCp9t3zEjwfX34o3ZoCjSYyNz+pjwpxJcjEiTryHEtZEfUR
s1XMrDu/NNyqvX+ujvv7A8FvmktiY+d8mnIxhzWtcoxmWIQNUDdDkd9FpahREf7N
Nop19ywg15gXP2fa21lZXtOBwT/vcm1uVIMG2sWW1WCJl+1LbPmfEADQSYij4A0f
liAErAoTvaZn6KktLzQYRo3kO8F/akVDt/fJlkTbIXxwMKhcw5h7ItsuCJHIOZhT
cYnsu6PJjWpvHfPxMB8WU7AIbwq9pz8oljKLJqYaABt7u7hGz8xcrxrWjTlWSLfv
MEbwCZP6PexUw3yKL1mtW4mGNpsA51BJTakXVm/30ePET8+uid52mTwXtSvEfT8l
B07IxQEvIVna8vEm6SZLj++g8Yy970ei3r/FD/4Duku/g/q1dmHtZxONGc80BNR9
knez3C/L1RbzGGnxZ/uI5IOwnzxVv9r7UYdQx2eMSz5kz0iTY1AnQdK40xFsd1hJ
c3dWTTKI/anKS9CyWKy7WmcImBK1fISc06cCsZwA0pxE4DTp1AsGAmBg5liaow6Y
7zqRipuPgZ+5ROVyelX8sCYJPU03wihMpzB5dxZ8DUQ49UGGHzSE5tiIt5+M/Tq4
0fhP+H3VPEv6Wn51hET4+09zTBcqL5wGYSWXKir2ygNUTNnm4uhBb2mgyA8tH6dE
2Gud6RkgIkTtcaBzBBx3OSVXnToioxeNGh0mjSsRuupinbJRlAkJnBAXvulosiIm
eLCfmersKiTPe4WWxUYbpJ9q1yVVZOvHrXMBrxdOlEreVvClnLWR6p5WkuWM3mUQ
DFLBEnWRVjuVYHlRnsu/9yf4X1vazxHyCtxvygkEnry55Yl3D3P+vHStOv36Qw15
PotmiSRISOzuIFkSRLC47i3cLtnKLkZ3BiyMrzpbO4sGNMPoXo/lErT7O4VFh2HR
H2FGti+zMX35LXUlg8nEMdms6mgKvgwIbN8KiVavZO7LkzCvJ6RXbCVu73Md4Pgq
z2aYrP4RxsT8V65FMjE6VI/4IIRqLarJl9OewkdR3mRnc9sd4tcPPVmPapqvX+LF
WaRQyFw0p3+HwKjkH66AuCXpuN6L4GdAtTtR85ZmzlYQ/04i5SGSHWf6rEdvyNNz
G6ZfBkSDtJ5gkpmywuCpJgA/4dJ9MoHpzKjrcczKF7nJKN/oHTuYU830pGN27mls
yaG6whyow6sNULSs/0ZwqIohlCWH1IwpRWT0ihBAcgcwP5nHJPOPQZkMH+/R7ZmC
x4zTm9x/YUic+UJVbNlKXkxQJjz2oxDDtGJbmaAGY/tluPwmQIILgRK1aajs9wSQ
r7YCBoFeUE+rxcXvLcWuASxtvnOqeJYrk3jg+17kp8j6JYnprmRWm7BLtH4o9tbf
TFKfBxGGFXsE5lu23mAWwlzQIdMhxb546pqxFXeZicA3cKZuuS+OPaYdutYqrcLr
wt+SFUblhMr6c0YAnv9T1kxiASlQlTn12X5NOtY4rRxBREHvkA+7DY6LiYSwJ5D0
rL9CzkGYQORoKliv9Gr/5k/f7pZXX8SvNwTv+GrCURKVK/TT1JX8ZGbWPRZRVPyZ
Fx1JpMGJMNj+YUh+jxaQhZ9jvi5LqBibZ7HRzRmNWQ65xLITMVrTMb2RmU0kI9Iu
kc/S6qv2fgizNnj9PuHlyLcr5doPx/5jGdLhu/jBTnTYhmxTCpZ7Avn8rLhxYO5P
f/P5OdTRiBOhTnKz/nYdhOh39B3SyBoycMARybAngEVH1nSmVS7VvPTqIl+vuaAB
9AwUMhxgKo7D7Q19WsCLgEEB2YZdStxnhuij/EEmtz00UsKTMAtIw2SY7iV6Z4k+
UpwTA3NlJ17ArgG2tyZJLE/+SS8gEHEtavICkOTlZ0y3BNwrE+WGvHVBTknvULbt
JLWJC8cHJkdt+MAvHvleuVm6coTu/3OnLthm1R3H/+ji4t+5Z46Nis7I5eNt2jOK
OcxJ0KOiVXvmEqRGnxmeEzIv4biw+GYowSyaDOyzom5RBzo/hNkK3at/kp+/BfBs
hoO2rYfdbP9T7rmxYec8LxbFwPdefOapOCLrTK5jtGtD2vOaSwLPhlaX5WSYuit1
0OFDVzZLUx2pDdt34PwG+ADRaC4nL3DDrW/eVHCx1ofcJDJQcTXlhXgYLGHDpgif
ZDm7Rs2M4norLXIC8+bOENjUKFgfmpEBUIX7pEvwYe5yAP2hjcJsRm2g/bz4Ah2r
NI9wfeDpF1s7rg8Aegm5IjLVpn/7PrgKruLxpx5R+TFJTf9a3wvyXrVRKvOMEJXy
ZnwopiOMXCzHZRBe5PvcBG6Cc9lDD6k30HbdYyuqcw5b8AOmT7xlqtQCk7si5Izr
YOU0K+wK++bZOHkkNa9rmijsbLYPMkbanT+Os7tjp2wAGYpyAmBCdsO62bCfxpis
ieToJcnKFzDbmF79EoYmrFDQuF64pSMXKxT8Tmj+azZb0eVaMdOFdqm/XLADMKph
sLeuyH7VhYbbEnlQkczuFt4eM+n6IUZpcdUw81h0YHrXVCJW1Gx0YfyniT6MmWAl
xj1YScul0Bm0sWlvuNpoWwCh4Un700PnGBUsU7CU3kKm/+0bf7Pe4YDd1+xKzWP1
JtYDiJjASxaGOdi8IOnp8gQyJl93aF/xDj9kJfaAZm2/f3YFZgdd0cBUlPBOtXnU
ykXkNFQeEZP+PYgXChuCQb9sxdafEU8Y7Ni+fs11Qsvf89inafTUGGQD4ZtiP2UB
IC2tq6KSbxmijdZzgDszNOp1QnXR9qUfMBSgcZdFbYgEqNQ0CDvIItMS012rqzCK
LzzmW2t+eRdM1xh0qlfFrfIxn9A25UjUYJwgZi/FIci23EqWK616uPJy9hWn0PGh
hrpKi6fHiykfO4m30b+AeWcbY+MCiLr/lc+bWzhbGeJV7tKZdybU5ZxYxV8pAYCo
zIQ1+OCvl4AzE2wZ1vuPUN8Nzxt0yhtV4AxSw74myW5pCkyvxsoFb6ty8h0zjKq9
3X8H7HmMQwh1BPO98x5Dy/xTUoW4t2Fjeoct0fuygZEsRKGPpXwvCQMDsFesZ8JJ
ElF7FC5/5838Vd/4zxjboG9V92dKE6CsFS12U3pcKrKgpGTUJarOCAPGsRD26FmE
2VyGaU0qjVKEX9de0mhv/uub0jnD979wE49hNylBpmLEk2Y2UtJy5JrUCaFNdI+E
wepA+FHyh1codC1NzHVt/lvyFNwo1F7Hz9GwCSdyLradAr1Q2KBptcBIDp7EsP9Q
DoBqYDc9oUE6GQwzF+++GDW1UMCoq/PH0A1weCeTlZnVuIS+DPkQkHGwixDppxZi
7aZuwssWw3LKIEHCwyA8XeSZe2VoBA59Sufl1WWpSPAzokl1uHK8bc6EzZ9E6+5b
IsHPTSZArU7k8QCvHBNEivU7V51cARBF2pxdTj2J7M2Jsr95lt2kT5q8KPMV7HRn
dL9Tf+tIgzI4aIQu+TPBj29QqlSLZiI40XR/wkvgfFtLunEhpwKVTwh82cWOfxyn
IsuNJmL/tm8qsB78OE38geoeonwtXhCoe/UBHIsggRSlkjMOuF4DF8GcvB+IR8rb
/xI4ZCRRLUIXZjIh/vOFE4qXCJFrWiu+2hcwuo8WbcxTKYD7VsB9H1y5KjeIe0BF
Ge+EF3DkQhfy4WnK5OJHSbcbQ+Y2wVJQrtmukp9KhYj+kPdzl4d+AVcnMfbyI7FL
Fs0rvcqXbPEJS0hfeLyTssdK5TFAuIH3LHSGM2idwKsSj+udeLuEdGgEuIuO+jrj
M4pSLfKEpTngjmsngdJUNzosbjwvVviQJBim9Mo4VJWGa5JUXp5THZsgCKImOSHJ
BfQiQDPxcqXT9Vt3JBzxroBM2CqDCCrCWVMnFgHBgtSTIX6aXQywwo2+Gl9rHhc5
UwDJljWq0n7t5N8IhEVikeY5lbp8TQ0z/SBtetAdJjWyiWeu2TomF+SpATSFMXZa
MIB3dKG9A3lAZlcB0s33oWbU/js8KrCystXgEJ6Bya0VsdmEsnqifJTLgBxqvCL5
QRqcvxBoQHEm9pviKTs0UT+hcHsqmMmd5XK1vGeCvpcItCVGzFW/M2+CMq6v2Wob
nK5dxq5lMZCgHnRUIJ7L6JUL+enA2nHgg+QVi5UC92nP2ZXt6+7hxbbAQTg/hkx1
qTCgjX7N5+jSLVFUkLVIbW8WuQJoPyFk6M67ZNKigVSiZD2DWcsH8OGMF2RLLx33
Gw9F+v/u9n6nBGblq55gdqDFML/Exm3xdN9xH/0UpWOU6Yto389zyWKLeBLVpiIU
MlB90slBMcWXlm0Y1XZwdCFIoWzqjFEnDuFTRXpdxcRAPQyhUrAqoAIDW7ZopBhA
Zr4U5a4E8XZs0hkhBYRmvIRGATLVrfRFu8AIWN+l16tZ9sqjvtncifDof407sywf
tAjRhBOdxgrcUdA1IY7o8NnsKPCS6jbzD2SRTWvql1SPrIjRURjtuao6yCEUh/WU
qkOcDjw2be9ODqUf1itYnUbLn+X4m/pvNNO5jwZo0rG1G32vINfKeBEHSTNdq6gE
LCjDcRfB7QY0zMpKz5TLtmHGyhZBgxbHAKqqdn/N402vZqyJ3dS8J2n1aGm3T568
iBAh5JkD5WcvxlyqGLp+eeh4hUvhgXBwZul4jVlMWw3KEWmt6vG4dSckcH0HTQYm
06cc/xsQYgQQ7gs/x3M7VgOny6QNh38LMJUpNNE+n09YJ1hxz/5KereenetdvXj4
WtULzOYLnbPps7raqQVkbKuAlzcynPOOPIGGGJpExkV18TCHVEMIVF747HkepWMi
oXllCpZkoES2anKlBY3tr6hUZXDfhcpeuJlMSqP8h8i7D9nBDdobvWdJpG6wks6z
Zj/7p5MR8QeAfsgwSNjoUssCsKcSjOlOrMf69Cmd2OwoxEJMnmYkQxk//c+iyrSS
IZk7WXZuSHkeHBVV40Jy4lP1I7bdBMc17HI/8eVOV3f2Eg4oLjnCtZJJa1HVA97W
NJYiwcHgGs43CaAbXG8ZqYDjQj4t1tuRmfkWFU1RFQPVhk6WHC17kKhrb3gqGuWw
ghFSZevnFiYnjSoVH0sF5ErFaMoVJGOnUJxGsp167QYfypHOMCYsbFRLy3gaMHjg
JqN059Dp5VS/mfvvDAsoXBW7eL9sjCSJOA4jXApkY0F64DPEb5VkLywoFKu87h4W
9tBvMIvTIGq1RkrGw0qv88r/4ho0L/iHjWwI3l/7Gbi7UtdyHo3Aoy/YQ7M45HV5
yjaZVCVEekxoDN0qaStO9evxSGVgV3DgyjV+HItjzpN4RpaLPu+DqNf/s+ejObbq
Dp7I5NjQy5R1fne7LIz4SmbC1l/hl51EA2NX3iK7+U5iUcXxXc3yx0SyjZgTL4QM
q0Hm8vkZo3DEYTT42lpnHR6uP05uSmGzJbIPDZDqoIyZWIu9jZmLPhuNzFGfFneb
FrSU4p1ps+ZgWAP8btnicNammvhrFrP0uf7WTYXx/uJ5Pv8MzoXF57u6PG+bIbHP
Cl1jpvGWOH8UbzuePgRWYQpiyS+ilwl8GSkl3n4kIMB9Ihn52n8nhFstJskqrRJW
4XGBGRzH1RmM1xkUE7Jk5bxN+ud5KXRaKdaa10nsDSWfFAVMP/E2ICl3SlOmM2Av
adqXyhs/MZxAc0weOG7Gm42EyQeN+6K9gnjIw2BWxvl2pfu+UueH7AEBj0aEXQ2b
/O+BdcH5RB2Zzaq6xiiwcotV1npx+YgSG59/1JFNJ1mdq6H2JP2o281tU/jzfmDy
cXKTZ4JWz+Pfu8sbnDRVGfVnMxa/hfheeoJIjR3rXFLDeDIbABKkdSeS7mJ40hvf
qZiO03qCknD9mANJmItj0QI1ep2BrYUzyTVv4xgL/Qt+eqTSQXMafzO3UkziVwD1
5aHXdx2Aw/qAKEAuuEvHwzL8G2XA2kuhjEHireDzL8xtKxdbljMxcH4XeKKfd3ay
QjrnOj/sMizKB8lC62JiQFvIvLK+vdPjYyIBmIH6eGx6HwKcgQKV6d9VY94IxxV0
uAaLRM0NgfT1eQeEBSzs0RR9MJaSbHc2RmepsFqH/j/LEIK4huc67eLjwGhKx8cM
3HmaE01Hy+zWRaPJLonD77TVWrIO61pEhCyAGBTfW9xeFX3TIfk3mqcwS+4kSnxZ
lEWQIWm/cX2r8dE6wZ1WkHmRGWsCMn8PRkLtPFV8oxeyxNQDQfYtSeKMi0Swr0L7
dWBPD91xj0Iu4h9dcpH03HQl9SydBPKPMk/911xElTYi1mHEtLAdz+6Wk3KdmPzX
pKsYkpOLW6BLttG0rAZPZ45a/w2aZ1E2M6vEuChCpZ/s6OuIrSvCVQTjVTu3Zib8
5cBIRVqqHVetYxfHpnaLma6F1vTsmubQJZT1w43XJS2FcWThTUp9I4ut9sjvjKVl
Wq8GHzmRaf2m0zPmyRE6np1alTVBzwxNfnc/euWlarfiDQdUZdI8lR+SLrvvgTES
Sqb6ByST9Ul+budadWyujGEIBq9ilMl6BYZ7GIowr20huKWFG0R+jYmJfv5/nWFQ
BbfOnrrEMjKtPb6Jo6EoZY1wo308Qkx7o/QIIZoEla0unABU+rrQ5GnMHyad0O1y
WFnfSOX9j5+bGPcKEXl8yaKusRmqA1kCrhkfg5mjHnmF12T7gKz2zbF5NxiciHQs
zgpRwl6cbc+WVHWuzM/lLtCABR4VmpyhPwVTYqe+J+0xXDWmZnW8EjaCwrnm6PLK
KtoQA2bTXcDRCscGX5MkexSdpDjf2+4W2XctBayWeNi1mkx61vV4Yicq2BI6AOle
cdrkMrxQdPGc5ndMl1Y/tSCJkoq96jpWMr3bzmEn9SP8mw7YJWqcFa/60YbptHRB
AxQOlSgFa8oC3h7tON3E0lhDXBfScXZlzbJbCM+zwfOV1zdZTlvGwWElTTu5s5/X
0NJlvrFp8T8hicVSSjVChqGtko2pOIRlsa4vlmfpdYeU3Qpwnfk45qZGE1RYes6m
ozYveQYvJdS0MSVl+myyEYFtztkKCvjPHkQKNW7nA0SY9MorSVlFfAHK5jnio/CA
VJmOWR3ALuqHLODr1kW+HvSmzV+08hFWJ1Cg0qzfFu3at8t1qlS6F0SJCZKEbPpN
M6A6Fc/W4/LK2l8JZNBEZt7fShSKJ+GXJ6uCy5B9xdqiO1PzaVVj6BPQRHMg2+Cl
vNswidf/ZMQWtUcvI3mgiWr+dq/62ZJOGaZaKoKAppVvMICXNueU+7/5GPIG4Pk0
yNx5v+EDvM6NNYP0h+IHkBRQa1oozwZPr1h19BIHbCLnWTXnIIARVKOx8pn6MW/p
1f0kxnfm5nDN+pcl5NdZRgpm8ByhQtU7xRsQ4T3E6uaPHSanQvlUon/cY2P/W7vB
3IimfyJfFUVVnKsjbGVoWJ0HsGHuUzDKVqPDfj9R4mcjhNObV4gkq96c5lMspIHy
wKjzuyfryhyDa6i8k7h5SnYj+k43TsoFLQl7zN4g3tWMv4uMFhE5X7ATjWX3ckwA
mH1yjS8+HrnptniGOD2Hp/66YLvR4Z5S/Hw58D6temxI2Fj7JlC/OUsWEQbO0Vef
xVTEpvW1a7f/3zrC/FImOCBuJnKYrIhjK8d33H8QbA8QLzAHdOGFrMVGZAcBXaFt
VZ1XoTxx2KTnO2DTwUVx3LuIXNR2PGpGqTC62mN0VN3biodz4mEAK4EtfbPVmqTL
0ENrE+sis6DsV7dYsNvcpFfCZSbeuEFiqr4UpVqjN9KqihB7gVhqqO4KvqbPS0ZR
GhOUmDLD16xnOGBzfH5nThmxJ/75CNcLCKcUfZa3IpLQWXATo2GSMOm/MfBjgI9B
/5xCU2bGYCFKOtyZpzrl/09IQuV58bybDhd5ve1z0s6W8nFX31W5APGMzEXJQM1R
H2vI/rGbfiKmXvsfp577damwVIMc4UjMO/qrFxqn5tzmtPlCBjqqllDWgvY1ggQA
7dsKCYXkMbafkeKzOlawprizyKN4SJo8/29blys9vcOg04fWcVu9nEh4qgX7pLVd
Z7qQZeviZonBsso+GvTuODJQiWNFIusFZsBhROmjbHQCLyvjizPQXoJJRF0EQft+
FFpeQlkSyevOfAljdTf5dad7bLPCjF7RBKT54yXKspzH4BFSScg0NkClhE66UV3L
MNDuw6N3hev2gdZsxlhtZ0nvE53UryUDdGbEPAXtBNoYGdBIcd6SRnnqVKLa6ZmP
/25WqZm5vm+r4Txw8oue/+DjxnRR8M6KOrCZxMSPVVpx0b8j1z+d7gOYt0MgZTxL
lSdHsZSaODZFV5ltxK3Sk6f1uSGY6XzM183nWOAWMU4yywtMtN6/iAG4iTVpLgJ6
tA0+3GsTYD24twE11J8VmIFqqY/RrprwnzTEKVJybKlBqnDaRvNTKsqv+aFSoBWJ
s+35mDGHv67NBPvNqU9iMU9L3DbTJgTtfGXvuh9CT3Ra1LdCjMlpkl+7tcXxknw3
4aADRNM59888pEmeoYiB4qycGmli4qQ7TUkZ8a/JH4JbqbzUYxS4RhzD8TRkGETD
JGk1deWd7S0MhrjPHclRvMuQ7io8ZoweA2s6QNTPGg/FRoF+ND/TR9LUh61Knwq5
18b+ZNae14Uu3Q8ncJOIMH/wh4T9O6Kp/JETBlvVDVB+2eop9tgLJGTdaMghNip1
eMhcFmTtbVG+ukIcaJvlaZF6GnodOuRe08gzgcKlcjVQf00pV6g9iTAHW+Cw6gqR
ElswgcDlCBezo1kzUWBUfTroX6owLoyyH6eZl2sXw5pQOI/KeqqQeija0eLmldf+
Z9+OWKzBswH9pVK6KC2HBlBBUp+Nw3yOOPJfhyPrtFx+yPxs9t+yVvDssLThUz5K
CjJJwD/vm7zq47VZmhzDXnOH260wTTIkhNsacuXUDb8Ygv3T64DK0yCwNLdmXPQD
kPdRlBYGS057kNamfY9oospdzgXjVK0XqDT6gauQv84COaZ22Wj7avSMpHCoTnUS
VDrfi/dP557gl2EQwfAEOnitBTOlEuE7H5icE6hv0BdfWvI04M13H7AmNu9POQ7n
8HuT3Yw9xVVl0RhsgSpZS7fKrUuCzcevMoaGlFeOIj4OlYRK8UtQyjcKAZH3Rlj0
qG9fuDR70xS7hEOw+glpbQNIJJaiA9cB0TFfqRxuxfjVBGSFh66h0qxQYngpiNBK
tTw3JEiPo2XdYXdlvnmmgtqO9vxh/vyFUZ65fCKKXTP/S+lXxAUAEojI4cObDrEy
24OAyyDSjl5qJTWbO5KguiZovDXILiIzvPWVsDr2k9W3+WU+j4cN7HNPz4jDRohE
+1MxSTX5pTKR6iUFfhXA7ndFVkLAJuA74tCzLr80u0WnIFFDokq1G/AzJk2c+5yQ
quDD8gXTcNyh72sQe3uniYq7WhRvw3+m2TK1sBlNSZJMh+/Xpr9NLl2FbJf2y0xK
XvN+YGABviGBcpVW/sDUfU1Xc6FfhrmwyOGF/Rjx3wOkQ0VQEaP2br0r7/v0yAJe
3hGcMvQWnCXhbM0tjfelwmjEXWpl9RQwfY4XQTvyDknDs33kvb95CmyLxTP2+5rP
tH95RSfZJbe/5wKBcYJy30qQLId+YyaxgcZGHkx7hZfAVXq8l7PAazX9xtCcg7Sd
YhwX+AE7HEYyUMJuCCJJpiSSHtzgV0WmIo0B1AiGbV8TRBVJRtUaXNR9dV5/sabr
dXudW+bvYIeJAz5gL/iMD7OCatrE0CUfVjlxor5WQ3CkMyFhKWBxqssTGrlrgQBN
G7Pjw5l6if1SgghenlPLmz5keD7fjDcUkA00IA02K8k7vaa4IRKbBUAa51IFAyNs
TDDZTA/lEGGn7ZWpi5BGU52mQMs0q0DMm04VYYRvrOiLeE/I4msLIT1VUDTD5O0s
KDJFjYlTtAXf8TaUk2etYXK38EL1gLF9b9v3/c/fX5inOEGkrVk0/TBVekjr52SK
3bWk3K1iLtP09SaaIIZ/wcLd2WylNvrTNP+yDB6W2kcAmE+FxusbX0XpGIW6xyOD
nUp0ZLKkjTkYIRKgbKyfbKmTVJIEDf/a/dnc/yMvmuC0ulUQvaZTDe8VD5YkN+md
TjI81AXtUpgZdClqHVDLXFK82BZX/6Mk2ciV75jbYL6Jx9YisOiXUV7hKL88towN
IL6yGnsnbW86DDlhXNPXfy2kZTf3VNGSQXcMomhX4zuxyR2AIqKN6RMVVtVWyVIX
PS9hoVQExBBNULqcJUoIG3NeZ/FCbuNJ5FRWSl7w3H2V/6MQel1fcqKR6uARkgZ7
FgxMEg+C/3VFAFiX3JsXrrJbRQb56EIcqdf3jnmOxcwE4Z6wBu2g56jP6G0lghWi
8WmDoizIrENTBWknGkd7NP8L/gXAz+v7sCFfP8UMSKOqh1IOWuHNDMZsUezcuC83
eqh7Gw+P1wTo8xIMNYuNhY3HMSJGAogAl5NlLCy2lkEYOPXotpt9LUlkJUdsTQRp
xSzE7B3ZnHe0LW8HtWlYCE8BMfdIX/EibzpvFVm/b5LFKlLkamg0+/AoVGS9tzr2
7rPCAxZH7ipcJOfTn8sSRKtLFeuj9yBxzpOjHZq3CjWZA2y2OMGvTCrbvc5zKgo7
DB4PBJhhEHPEqs4BQPoQpfM9o5HWaoIAJbprLA1NqXf49g9G9l6+ecwpjMHq5uh0
S8Y6dHTKAfT2BfODFXkuwdGGrnw3skbObytm//REMPV21F/Wx30eSXwTB6yuRElx
Zgg8idDS6KWdQ2TMbTNu+XshKx0eiGX6uXBFmL7XD8UwLcjv4pqL0N6lPzoVrqUD
npzJ5RYKici7Do7R74Rbqa47aKABVCmxfDXAUQGygg+GS11IAaeKrQMneHy5C5lF
+gcLbIm26nHRWPXFIy5GTq2ZH4JgwpSFz4dENormp2UH70N7ZRKLN+3kJZFcQyhl
hCxwVi4wwkuqpjmXYPt7v7GDr7VRZTLmaUIX1efdeFoU3R7S/gPYrwkKrLiDvGoy
q3Mgv501d4ZNLfucyHTaSOMB/nr/K6sdDGZ/vXpgyMESZB4c/qKH6i6yjTuyRmlo
J2A8nMJSL6mRPnkDjB0hZ8e3syxMXsAIxtnChmTMCcKIIPT2m1DooTIQddn2LIWh
E9xlQikIIIZKPfaEnj4E1v3NM/0sjSUcBrhUjzGufllYeuP6mXbEGZpdkDmlhGVt
9udwzCPlLQTRQc3LG4ZLzqvK+xMGyflptCs10RNPEcjKzwR9mdCYNey49vmFl6p7
GnbS2vq3zN+ZSXB5sptz+wrHp0ftoRjEMi0sKUCHyStS0+6AaEGJ7S3ZOIVn5pHG
5bZRvylm/uSDhoawDVjmzo+eTjK4pJfSOlqlSfXVrHM9MUXLLbH/oq6dmmZaCm33
lveeDuUeubVPE43RqqDUW9TEPmw8PeCedDpBS2JOfbGluRZ/x9GjUL8SC0ZY4glA
bBXF0tmpaIdtquXUZWMwDU65Ap9KtgNTYurGJSu+wRcRxw37IAN7lWERkpnnUc3S
61Fi/OMpB9E5iJBvNWQepLgyikXlctuLH/7lVjY8KEfJAaI7be/rqIcVfOHBPHtB
HdDwgED9dqbak3FybFLSyNbmj/jsp3mgPVPTuAap+7XK5qvj55x2l9lsefxjF97r
Gn6UOxxT4ryjCgMAuw3durg+LttXD28oNtuE/jLr+cBpfXs4QEpfAy95OnLHzKgo
M+Xfsqo/+7CtR/7O/ymim0qragwygObTN2WTJ3pzpAxw864ZJ8sgAA57KBUQNZR5
UNmujpw/U1QVh0phe+ArqG1zD+YrZsa0lGrcHqYjaT0nyRrG58amMMHPW9c5ilQM
rGDBOQc4wSByAZ++gt/fpR1C5pPqmnwUZkWqMwD1SUAVzX/fxJdbgM7XuyxO8flY
9IS/IeBWqiDEfBzk2jga/RaZtpIAceLWAo03l/TiMNQA3u2/r+abpXQhG0CMV3f3
rUY+Cg0P8zU53tl11WrTeKfasM+BnduwDYw3tI9vfU9soWLDSiQbFSFD0wC387+A
hdmKAGfcRYaDPElCdfLa04aeusoiPO2fqujk3tRUc9Qo7+t+D4dGqRpnCCKYzbMS
ZnQX8ugX/+MoPjRzTl5kp7VUHxLhCjSxYK9Gam7DZICPqTq5CVJvbvGb2ccH0Zg7
Vr1t8LyS15/+9w0kJfIL72yY0u0C6jQOHq1bqNCWZLlR369WX2QhB/N6I5NGx3To
q1OuHOMoTJTdr49qpVXgEvzotDTleSKMcWvij+lnFn1s/Tvb5Uof12+Es1jotDqR
+z4g7Q+s+HMInQhlDXL7IFozB4XoRA0RalrON0RhzU119f3vdt81HysLZ4nyNgNq
U8nQgE0mgHiKLEgPBPPAFM4bEBFdB53vHUffilnOEKghsobfe1QVuBo++FS/9vTU
rSFR0sp/ytB92qEzFn+2ueEIsYLm7NxkTbZrEG5aIBmipfqib+qSZ/+b7L9g4eYz
sjisiskbuRfKOyLg3fMJFaSqTphM3lQzroh6eDmZ6h9GgI8nyve0yofXOBtS2dao
SbRKiDSRgI2THqAjjPoR1fZlBmHfVb7IX7Of+ZnKW5jrX80m7f3iwU53fLQy1UiA
eD3ToTNN+j+q71qwToiBJ9KvlUbUAd++Pno4/5Z6uG4XWrtwxQS/d3XG/WDF7Su6
ydEJ+KDc1VpfX/CaIVC3V2Xih/GkaJGRgzVseF5GEPu8f8MQuB3vagK8R/VwAEej
5SRt1d4j7V8lBSPsiAXDhpZBRD0LfAil2r9gYiZWiEZx7kt5vvVhedSDuKrOSSz9
HPnTT0jJeX2sOUo9MuxI+f7Gt3ZGQZuUrHKHsmMIfTuxCH9ojclK2HtsLqZfsIJy
pJV2pOWeIS5FzDnV7t4g8z2xvrhbP2kuk9zfUusBaqxQQ/baQbdgQVDXE6OQRcZN
tuD/d2+h/39IcDuJmWi51rusXDYISe8+3nC3DLS+J7k6lPjqlkDMXj21ZVv8kgsS
BM8ZVjcIZ3eAnYKRGonoRELvFL0qtxVD53KcP+zX2nAoJSIWYKiTKiAy5ZQ0XZll
lPHdikWuettBzYi2N9cavrkds6hbYIpw0fb8h3zB3G87Xq1ASzRkLJwBv8t0hmx/
uz4ipUDUMjAGgNa3/m6gWkXgFDgZjVWOf+bvDX4mM3oC48020ZIDgLqGl+bxtkLs
MO35yYaOn4K72gQJcl+YgtkC0RsGM1+HMsUh/e/8kxSvoqFTaHTTqMZbpnjAUK1a
iZkBs3r627tuMQbOXHtmbtAHuOoBfWDT+EkMZVypgM2s0C8jHVqKNZN11LvskB9e
U6Ds5awX2E26aNLSbaIaMuhHmj1WGDjrvdsgvt8itHkRrgSytlzb8dVBpZWP4sdy
QseBssHnlfJHnQXgnCCDsrcBzhmbpgK4ZUYQa3N0WpkFQ0WVEFDHXKNp62gyQ0U0
y0NuiI6e/Q7pfC+mwBxl8hzTn01e4AOtTxuXnHPYMdhEzVj8fcScUEJzVowohUFZ
baOCrgrNdGHoS1Wjm28FFajcSP31IKxJD6IeYh6rs+ShZea4MqxVvOolPx8ochZ/
prjHN966p4XIc6EkImc8VHCRmfz9cNbaiuyo13r2FLX+pD7jfIV4qcSt6upqMW3f
047R1NpWqIBQV793MAqXv82V2ouXwGVbYDnShEOY06UeloFXtfaTR4isvwgW9t+f
mtZ4HYXqOpC568ssxQy2oOLT2kMomancpKAytnw3kQ+mtH1xKdDsR6Di3eja1WRO
wwCjF+0DYnrP+iijXV3hQmqjg2No43qES1aybiVfj8knIczK87T5dKh7rBs6O88R
6/pc+BPhTpXOq/y6CCoqe+KO7mQJnpqtCkFHoKcgXwWF2oMv++GQn42OaiemEoO5
Rid7mPvBW/pPVS4M011QWM3zORDej7B00ZXt6UPWC/QKg4HTb3XGOTRGKFl4SP3H
ZfAqCShi5OK+9Hc7LxOAhyWsM25hH794+WxXZsGQQEf2FuSpH8fiqD3f+EsshNum
SFknAS1pfHbLOJxOIEkDURQFjlQGf0DGWhhWqeG0C11B60azZrA4fBHsqXxPvqUi
BRlZr6eyzhgxHYcJL/9NQ5K0jeDxz61+cWyxAZK1TilMEfGrirdlnulJYWc6eIkh
oXhmGWVRoozs6aISeIvPkuAlEaTWPT783jp4Fp2e202me6s6AgFcHaOsYVcInD1q
lvg+R2Mk6t4vV0L8q7kLj0MbjFDQ1X+NwTjxj3PvXi8QUX/F4xA4ndZBUCtqrqka
6UVtLLB0dBPlbJA5di1IIHm/sDNoZ9DI8SQd92dx7ksWYkBJLHRYugGiLH1fLp3F
liTANL6ioFxCfBEE6qKt1K5iiY3wuM9an5y67wSmR4TJUaqRela7Hqh8TuZSxyur
+Z8yZ9o9WgxyYTKFLqtk/lc292uQT1phQu9kc69e0+6PkNKkFqUoXM6/XLi9257a
HzzbXnszrNqKseUSgXzU4e4dOpTeWOwo+hmxC4tpvG+su4dvenQXU6cqUMCbQpE4
23kEG7oaDB5hrSd1qOELXgsI81YC3saniCVxD4UB1Idn2xPbAYZXkbDPhJrfmvtn
uE/WM5OjaTQgznVUUDBKpUp2xnF3rAC8sgLyCvzI87wgh/mB+xhOHOL8lxqPJGaf
/pO0zcp3kGpvyr2yNLWGQfwA5AHzois0suUgZy9PDtXDSWZHXLkdqDf17b+wE63y
eeqnzkGIAaBm39scgkAQg5JFulCSm7Q8UQvKt92s0wRJ+8IqAvezuZbpg0/y5IRq
Pyp76RVd8izcU9pMh9YmryabLXfqVyZflN5CZaZsqyZCUT06AkpImEaw3wl7exM0
LlM4L8O1rsn0JwtCiNO/DqZwOCA753AoBGd0Wjc78q46rmBMx2ttFKMgNoQOJdNF
Uponpk8IA7aChHr3ddWBfQ8lQqARNckUAgQlQLJyuT+FCS+HP3Wz1GSTmazaAG39
du5QKCMrSDktF8yygiZrwkV05bAzFu/1bXwTFBT2x7m0ir7jjbRWSL+bviGzOT5b
OI7rJpSndb/y866ScfbVkD0S0LSLDWa/PrPZCSCKWEx42elYM0F0K5OYcy2aZEYM
4CaTsW9n/Sf0yzFCsZCjF034sFcjQHaOn2Aul9XbAO/NRdnnopUArOQlhz0whLjs
dK+AvlF3v5aNfiBAMAOcnGHYqkihEtPEmb9gR0s9WXh42DFuyT3u4UhHYMOL4JHW
ULZ7N2ifUOsAI/G1l0EWEU+JP/fYa5utlU5dhIAGE8xjay2oWrVMzwCSFSpKFMDf
Y3OfT7lXSU3BNNN2Mx94ZXNOvDmUMcCzLeo8S/rw8lLqXiDJOCJpozaClq1D6rSz
RcwZjvhy1IR0DXzxeoS93XRFgOMOyMmz9AewFLVox6rsdcy62Ch9Qy+pzEkFvgov
gl42ww4Hm2MwhgNGPC46LZwPRZcelhKZY9tmTRWPi48rvBMDVcf3kemoq3XFmxOD
Wo1U6QmzdyU9Qic84ev28igCj+Ahs3EmLsRIwONItmmrccFCcI2bt7doj/U9OCGT
hDW6As5FD4fk7TkupZKhkzVNB8rhCEXsIef0Ow8svrCMAwMwZqjAphCTQiaAOYWe
RRvdRz/QASMcMazybZ44vwMCO/i25x1YWQO4TPR5iEQPftmA3QoBR12kTmTnxV8f
/cJkWUNmOZtkLrI6WBT3bu2tsIGkkdsRsuBQ6EZ9xL4TqIQYqQXWXfYLS2TLBnaf
SjeLT1GSDUmZypLhvHWS8LN3xLubQsEgCOhTK1jlNwEPKL/9roE+ExeaL9/OuUtv
obNZO9KBrkR/DMo/KprHhJhF9K2ZBmKi4hYBCfmosuer9rq8mT5GV7Dj8M+xlnvp
9/15iDrYfRjwWVL6w+NSjdhltfg91vGnSlXJ15bwLdV12/oe/86aWjuJM1PtNbiK
PzA2g4//BqWSPgNjuaadHlnAYNweK+sMzgg7mx6aVWZ3OIdo7B8L2Ve1aiDK6C44
9lb59f8WQ20vb6h0r1YRYLM47Spzz8ljnwarykpIK2xXn+GSez9zoCFCFU7ZUA2/
Sx/dLgUD1LVF2xQG/q+KYxGUAFYzijx8hU0LfrWfKJOEECGI6kLusPGyuec2U8wX
YdUdpIVBeHU9VYBAn90s5q/HKrrCiaf5hQVAwuxUFJApCQU2gwYSLE9yjgFlZLW+
inGnTbfP9+OfDxWs+qaJUF+EofpBolpgyt1v1TksX4g=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TKax6/9OItUAVr0VlXs65FOxAmEJIFn5deEEykqv6E7zDCos522mxcqwAW58kdy3
NcVqrmpa/mnTMgcmaR+o/CCSbxLQHp4IuXHW80oONQOYMi4jlcDFkS3YFcZenS4f
H2t5/YrG2DbLt2Lj/V2/MDVYsaRtnfpCE4MsAVXYVmKZEBeyJAWqErw07U7ck10W
D90Danx6ljumaHxWzQcnkGwuZubjXEPO5lvQqNmWgpiJtEJsnh7U+OEsaIpFbQ9Z
RCvTXuh3P6SW7BTNhVxewEV+9poTZHi1X6YZrN2DQbq8K9DbDRgbBW6GZg7p4jjB
O+8iT4/SHJi8vSmawOZUyg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8800 )
`pragma protect data_block
UjWjy5WGWOv0bpGt5EJcg5w3Kt+RgZ/fhIsApJvJFEowV8RtmBhG7f1SB+lAOjAi
TU8IwcR7u0ogrBze6yn9t7A/3Zj22QwaGdzhqeYCuwt/a8tCqLbWKyP4fzLUbT+p
QclSKTeIR+vrnLpcu4kTTxCEognaA9AMIqwoJGl1jq36XkqIsMkpuR2XUf79du1n
UyO7VRleAeGsTkRka+HvkZRDRZKCd7qIPezVAzAIcCRHeCt/ckh4yTl4upIBPsJF
W7epyUUF4NC3kHc8c+3aTFa37mN1xZE6xbTlHnfLtzeL/NcNeTfLvIhpMPJBz1QX
2ODjY7UGsnHTPLyPzvKmMrrS+EqFusIZInNb2TvGLtifFAwaqJb3ilhaf3SJjUGT
8BV4eQCnecLvBNnKqbFg2YVL4p628pgh0oRYNC9BDTpoi2t0P5MWuZyJ8jH7jAZK
B9jzL34T/yVoRyOiTEsVQPmxJY+ZwR7y1RUsK2nEEbjQmZOZVbY0df+p5tQ+IU8k
6zjcEUyqm4cy0zeqEochTQ0tp14ro9wlA3BFp1EWiZXRVNwDlc4LfoOa4KoRWm6i
Oc70FcXk7tWrjwlp/bFcRL9prK/in37QmH6SnnKR3xbnGWK6EhrpfiW36p5Adh2a
2clmWfRpKyHPqoM6D3Uq2GjCl4Usn8Dx+V0EkuA/tRu5RLIJ8VhC6OEfF2gQpDQX
8n3i4L8KiI7LTVkcCXWcPVNncVF6rkgjYUx9m8OM2+YyykUXijwO2sZQAIiC6M0C
rEG/kEQF4JE9NbhC755Dk+Qo+s6eW/GpeG83vlIQLknIv2YizgtBYFCkoNnybBDT
a0wjRBa3Ukm77iuUQcTp0Js7QJrDQVRoHzwkqT6C2reVEqtQ6oMp6Y0gBwVElIo7
m7YD3rx24FVZE/lrO0vq9zZ6DHF4k7veiyClUV8QOMKMZ7J82vVCpbNbJMJSJcYu
7QN+z3A9+WYu81grNGrdYq4UvpB5khvlVvINh2l/bvBe58hmirBsgqY78sT8BHPq
CBE/1BffPj4hdD64sozvyJo8m0x4PUuFtQyvLCQTNkgZ+d4Fasd6BGBEm467HYmd
bWVCJ6JIzzdHHl/tSI2Lp02w+++hQv8VV0zjp6jK3FwvMCl0OSb6Ra6Y4Ox14FTP
I3mRm6WMYEkSba/gty7vWdD+Cy2krUJ0Gtv9HF1rx2b29qkfcBPdy0xc00sCnYQl
YPYedL5EenQwNja5LewRIkQoJwYTpeaioormfIgPo9gVlrMUazZBdPJX6HzK/n4V
f2Sw/wesOlf+ylLxsHZs/c7hU/dMQx+/bdNAKIDKxxOQ1EuMx6qdUIOND4N+Grtm
KcLxmXpKVzjvkr0xC/MZnWcHgIZIusZrkCAgK7xPfGIUF5SRbDArAsX3w92AHf2d
dXjmAfULXYVN3xxgY9XQHOTrh0muYEuHZJY5hd0U8m8YcZzEAfLeJmbrI22zrXTj
haXDx5t3AMXEO9lGjJ0Ewb+JjaTWSzg0OatfpFdqfi8FmQJYnKCHZsh3L2ow0Bf+
lmDsEx6D6N9wdiPmiba78oWOTWG0uNwhclrw72qU2hzDz2rQCgTMRT6lJXMdhMnx
TW0JC0PVV4Asy6a5aSaJZo9iuj74LGD/w2SjARDTSPf2PyiqVY5hYKR64q9i2Qwb
bH6tkGGFYLFg+zsGjWvARw3deEN4LXOOBU2pCeHKA/DMeLD2JADb/HAXmV2AEkxg
dCmgtpT/6qeMdM6pObk30vJzPhzeTlDaQk+k7X+2Ni1hklf2JizYp9vgpIZfkZsF
TLh2m6zB7xVE92WA61BXFmLX8qrDMRn/V8r15J26I4vljC9rMyJc1JFou1DwcZll
LcQdX8GkRkcTjssbLZlBSnWk7+ILHzRJ1FRN8p7+7qRP1djQu6d1UiFdEdhglonS
mpWEFgr9MrdGosi29w+buUBqQfsIsoxY8sKMciViOehZv0Sdhiw/ZlsXjY99/MCM
KhT3vGzGfPOTkfWjRywwgoz10bnIg+qSI3fGlTe5uSkXb3DTlAyMtex+IYvbFe6D
BGMHfKSIvxeUzFmCki5tgLw0dsPMoBpNLHfRfEYa9+ciVPRgI159WsuzvizbhO19
w+Jp3LM5aWLNzPZ/Ln3WDpACh/ieLTfS7tEYADqLudvW9icBlqwa5dVyfDDEMuQ/
MvoOto5o5facRpppYXRu8i/6vG2pxitmtZ4zj1hN7m7BSkiqGIPLHXHYVydFWSnp
Zn4aQZznH6jNONEMjgBMm16qtxFPzc7dUgMLN31m82ONtOkQOpL9cfpQWqq941T/
b7YAig22xs7YvRwzrW01KWt3YNqBQvjx8z5yonml5OeykXc/0kq0ryIKYGdBUnXO
VdohxT8I3UBgwrzJgyS7G7JLPwSxE9bEifBR8lfI0ZqDk83TXGweiZuGDvZayIvW
JyEKlgaGXgsGTsuiqljei3FY0iG98/AZjeToL3xLNWqI5bDFR7o+cpIaedcdKgV1
B3z02bZ8o+FmaA6HzUWmv297K4eogo+40iw69h8k2bs7g3+x3XFyZ/HCdBzDy6n4
G3Y1CM89M9fVxU+PCCszumlAGYHAN6f9hfTCf4dalVoC5z1ikARYEGHgzKTYrEqZ
eoScLPky2n7zP+RFNCZY9a4kp1EZTPPAMxqczuvPIcz5uvIzEZgCwySTGgo/0lGl
rWZbb6d5qbCyM3vBsT/axlSezuxKGTq16yk6vhClFXCXB4UOta1Ph/urOKS+1WIB
6zf1IJgn8fBGfe5PBvHoiymoA2Impot0grzeGp/Upu4L9IaOJx9YGz92v96vIyOl
g57YgKqxkN5dSOEQFuHDtlPFKi85fhzHH+8Mwj9PhRodqvn/z1+juJAlMjf5QyET
t9K/aYFmbdv6dBf1iTDzFsH2U401WBN642hps2plC67ea95Vd3rjXnpvS+NmxjHU
rNwIYFNKwJeD36x7TaLvW/RN9cOZDAL7UQ3m1Q9ONjk2jPpr4nAHkpW5SaNEP0+a
1e4qTWY/zo4yuYZnobtr0AfTqgwJKihNbJA/xmzn6rD715e/m+tkK6XMXtaBUjU2
wrMhzIdGVwZrrx0zVUgK0+S4o/S9EkajsT/4zn+1X41Xo+CDEyK18ptHOkd1OZBT
n3fJwzePxsSH/Ns1wzGBaiPCJ+/JKalbVCtqIbdR9UmpJAmUqse1iVelh/X7x90x
cFUMno8TAkWSwl5RD4J/9WAAEvhFUZWo9ZKqgzhYEE0TIFsVV+TzMZSl9WKJiNJm
TiE/X+vNjK9ESr6ZzfRXc6MVUDt+JdPF8NkairkKuqxb+uh/NacUSb45tU0VuIAP
7m2g5epU8rx7SolMrUgYjn+i40w2vuYosTtyE2IYumUmhGRsQnGhdmZaLLPC23eo
NOoAs1gm8SBba17b2ZV3Nwvey17cvqT8bakFQMxkdgk+L9MpVWIguoIOf87N7uBU
ZW4ArrupOsr5uLXeEoWpdNFipX30auL6osVxISuitbc+5nAyoksvbQSirRdDbOQS
9q02WovzIkApgoCamb2nf0gPeCOexp6nWoDc7YtIc7KVJdjhl2UJyGRK0ISW+vLR
1XTKfNnGCteMGB50pQMGLptpw1zXbk3AuZ5rzhXF95/bAYy77gyGjkE8E/2tUAIU
RS674vHGlhS8zUF/MOFmN2ENPLtQfGCvW91W3v0ZnqqzoM8RltOuId0zh0rf33kw
nQkmVdy39DWv1PKNZwyTIeUkTa2jhA8hkhbZB1MquP5/QUiZyKuMRZGhll7zVr3x
Soq7OTUsNtz2aI+Y/XI0rwbwDAdiDEbLjIfs0vwRcrZvNWy8Rx7PIpHVhFoOs019
ilblFvExCvztM8S68ow1nQYmsNA3t1JLK1KdoOHhUfyzAJ2jMmkY8Fg7q5ZaJK9P
a/aZBcGsw5C7vpzbdZmfO/R/ZxkjVdfhEGTwXqLYngyhsdyZwbnyWtRhULMpNNlp
E96TFI9Hf4xmxc78HS94VlHD/jayFccJUk/GoboZKGOtVOQsT+XNibOJhGz+KErN
dPtv7EzUP6qx14hHH73YCJK4rsM5ZljrMLRMPfoKYask1lmtN0acTbuRPKu/3oiy
YLN+12ojiohmdFnaXhxiOIH9G/dgKB0n6lcXrQci8n5TzFms8VfcDlOjlMRmtshP
ckANnxCOgfNzijyO2q/A/EsH6DEuVQGX/cn5Bx5IIRVp8nP3B5gKAZp2JE76Ctx1
jLigcxxQy+Jw00RzAmjuFAfdi3cpXVBxBEn7fkK9EooAYFEcU7cbhGLQEC/PJTmL
7w6n8HxlKkSLj2AFT2lgLuqcy3gBGaABVsGRbXXiROc9QdwMbY/twOt/WEqz+p/V
s+2h5eBzwP94ZoLa79OrlKo+Fx89oNXZ976suMFwQYrSPd7sUAMfK12c7WvW4E/i
gXpx+bWBBoUDWqFHo5+93rUFdTo3zsboW4Ph8dQLvi3E1DZ/io6Vu2f8cNKHSqv+
Yekzo++6UBbDivB8UEqltEjTbvlWowNBraaidWesT+xHV4Pdaf4pacgvv5BLMlP8
ur6zkkEWtcv7BMQWnoivr8Iq7f5msa2aDjGxMyv4DMKYjuwdZf4fxvi3B0PG+R92
3ijdt+mepEKrfo+TJpEQjyWz7d+FeSCKH6+oSY2fIu/xxEprgh8Vu4wSW/SLGOLu
3RprbRz5nyhj11J+nVFT1HFh0o1zk7qWAoFEzCtcGnNOlzuzu2UnudaB+V4kkj+q
URXviVrcbh3oOdh6jfvZK2he92cNslMOf/hG7Pfpjc3WDSoArbE1ukUOvlSR7Qkm
qrtNtC4wWVkbl14mM2bLOvcmRcqhEIALKZk9wm/xR+obEx8hyDFv31qPQZv6HKy0
XK38eyWqcuGx0IYqBsKziQh3DyYi3MVspWhj7+AvuzeamdRaMHqupvIHfFxnMI3v
tYhEVQCMwGuUSCjZw2JtQ41vLn8GxAeLCFX0ot8gRpbC+c4zkT2CBrQeJDPMen2O
rgWJVS29RUd1zcuuL8QA053Jgr4M28jzAcSFHkzdHGBNZeurHqitOV18YQ3pAhln
+H3CkYCv72WPzD5xdenlrKhTcoIDy3QT4K/HXNmfJbL+7wljvhiZC1Y9fakUh+lP
eDzCcLuFG5X4gbJfqC9v6xqNknD5JcONi8Ydu1lr+42VECdQoPIaOcqZxnAPNLfT
MigJ3M2F4Lx2PCSt/BWEzkAW9xH3Rq/FEPET9LlbK0tupQW6eeF649uZHb2/DnxE
aACqfgtwosEfNrKVv/9hneJRhxa5M4GOE6hAGMQ0gZicp5RYtRQ+60jad/tbKTMj
utrUYlF/iEG7o+VqyVe/WeuBmTpQoBHdYwgdxpFGOdfmdLGoagRIL3ZL48X7V/i6
UWHTU3pgxMsmkmRbNrK2gBhSsAoZEJxOEI26hJsyWSYNPklYTURfbHSTnFq+FQDK
wTvw2m4fEQPRX2KnQFwo/SBwXc/7kJ4RqjqFispZ+eGNQTfRwJ/SIl0EELHRon0j
4NhIXqPVESPXcrVBIN3Kllg8JB2U7VeJPMzHDYMQ1caBZOo/Y91yYcSE/1q+1HsB
RuztIyLe8nw9SttWvcq9K9Tfs47aC6jMCpcQMjgRH5NsRlrzIOmv+ib5si7v+li2
D0usHt37BPc+nDgyXVL2T40AwjtJ7w7Mgu4smVPokOJBCagWuQG6RusA7d6R/qz2
2B/bhKJFZtZAsD4zneXntaMPcamRba5Wce8JuzPQOeWcIF5sTi38Unswf7NtkX1R
2shjTEBbrNMgtT6n250a08g9Nlz6TxbgNzVpiZ65LdGOfKTTYfIvqK8LrNGdQNxy
CLJiZzpbXAhqQ/UGLguRTUPc/v/jjOlWAEagRmvJivy+8LzVt65cVPa1CWfVA8WG
vZw9wbRNXedMi/ALXj6Pb3WxqYSdjLRyoXs7veRzwR36CNRtEMhGlLRDdylN0I06
ctpSpUm4ShFwcS8NTipxapKDRdgYPDJqyt/E3YKhI9Lw7f5mycIxKwG8+comK66V
0ofN4D9DcmEGyhEA7WcBHUhu1Zc20gr8Hml/1/IEGXeJsE/91QP1ehka0f+guA60
f8ou4/xJm6psSEieH0xO09sJBPcFI2J9QaBfNIoFV7RsTbFwZMIMSm6pCYj/7zhN
YGChlRPlUkRl3eU2ph7s69xyfpP6hjfbdqaNjdHt8Dp7zftM1saCDZiA824q+0zA
jzd6uoN9+4e+gbFdIMeY2qfZlVM9yT/JireL9utqrXNKyJd1J6uuEJYOr9TQ3ElS
1+ihQl/qTnkFbHaf/4xWP9axBP4KBZAC7KfO2/wZF2zhCkAHHJX2RMnk8X0BOgKR
bY8378+zehwtkFvhWyl295l2jyHEpfeSqxEVpUbpAwSmhwnXRjkuKXfZWLvfilr4
L8ZbMWxYrf91HBr6jSjId5GKxzYun1xRyt2aAdlrQNIsPUBUeXiCwAF2ivxS2rQ8
kP6D9Q2VhhkAvXHxMTRkrfjC7hV4wo7pGN/WCucHbXFGzfO86oQCytcqYSQ2nUsU
Oo1GVmFWta02rR+IVTcsu1LoT8NOGUa+O+rsSYeAyS/8PP0nRQ+EScA+GZKMo5zq
gbDoZiI72Ei0PAPNtnC4STrshFIykm4a268fCkwNb9aY0YDxgpCb/8WeH9QME5Ff
tLsRRxCylZEBGfmt5hj+yQsq/cduYghtLXgNBtUZywohBR0MPsdMIU7SDK4n0me5
ownDZNMI+JHFMYE8X07RCHlk5jShdNGDNj40dOKf8w8Pu8y2gL2J2yaDLodmne+o
zxaOs7bYYRl9kpu/EoDo2DrJcgSE/yf3g/L58mrMFwA1AirOR6j2azdlgMNcZ1s1
93pfaUBxk1foNlGHrjR2zWB+cZTr82y1B8T0xBZF4CoYOl6Ti3/uVgX+PhvXylCl
KbcplikbNjdfam2KWbttJ6S4wDBpSWBL+6zWfdMQXIDI73gRkPxAQXk0kyYU36ea
6HaXjRBzkNBOwlsUZv+fcjUMaSpoX8GJb5bKFXQ8pzH16J5lHGfHt6Su6sRIPi6e
O3bSgeO4PZ0eY7lb+MaiiJa6uUWZEGvxLvdc9xKHT3RMYfTrI5Lv9xNOlFHr6diw
CGKkFOAhHLSZjEh469jVWuj3Q+2nFiJOgQi6RxSxY2MvSO5OmJMtvMFPWme0s3ey
L3B1gmKjtebwmq97Qla6QX2I7ZhWp3z2r0/X2qb+rWEwdkTRaMg/S09RdkktaTlN
dwV5+KPv1Jf+NeMvJryLIlx2uiRDJTpw/TcdYkUdREyCBSPJMvBG6M+ju8BzBYEg
7WkMYuJS1cEZCHIphpLvk6l+POmjMUgVPA7w/0ThLZvpdZn4PEMGvJISItFtgao8
3bUZb3mfGU3b0NW0kXuLeGXHifoA7b8i4LXqxXMgkuTrAreJmhivwbFkRDh8NTQj
CRimBQyASnsv4+S5m4jsuxmKQ5wS7p0tdNqiewAwTJfgSaXqKRUTJFE1+1Msgfwa
nzv2QsyxNF+7A3nz4RO7a66/tS1VaDzPZmCC4xGuP7IYemR7Zv7FzB5METMTlzch
0Omvu2eQbXmovRyWD01NlaDunwBvkdvy7mM0aQ6bhnLdx3vzZDI3GhvCvvQaixXK
1GBq5n4LOsXxpg6plV35kdi0ePDkP8oY03R5JkVLMtvnQrvbmbY5frPNkR78kC1D
d+pTv9vPai76flk4XV6aU2W7W7D/iXo3z9W51iI/qqS3lL/4vZe+zRhh8hsSzLgR
f+RK1SS1tNq9fJJVZXPc6VFWRKx8foAqXKexW9fr2QpaPRTKYmOvY60266qqssyM
ng1j1AdXRFSMJBcnkY8tgTGePaRVGM0+OhgpfUvTDS6UfEUhNHOM84hAXXm1dx/l
pUi3Pi73AdLj7gT3cX0QLtkvYq4KMETdb5LX6+QLTI0dkMEgh7M8sW97s0tB/jUd
Xj//CNHVTGeQud6IMZLX9R2Kc4RmvjEtralv4bKc7oD5tbNThpKErKqClys+elsW
54Xknov9/8djJuy/tI2OQi9yekelHAEHCNjs+J0z/cV7Q/4KnmvNbInKLkkksgew
Yq287Rba76VFV6pWMIks0M7ywgeZI93cK0+d+KNOiTJDM20uMYKBoy3gadavhVLb
oUgKcn6QoSiDLZ2Ei3go7dpKGpl/EK9DrMQDXWy8NOo5Yky9BcH6g5K7aLmOAQUT
IXDSo+va5thIPgzBNh+jK0O0gWSST3YtKKu8pPtCKVUgli4w/HA9Tzwx0UuBivBi
uc13jxSazPQH53ZEyjpiiHb1SDFmZLOCJC5fJIhIUtRfwypI++oJOaCyJfbcNkoC
H/RZuOFhCG/VMVc0z8rE/QEdLYX0lVNFC7nhQyDbtcUWxHyh5QDfHGyno+Gfn5lX
2cD3YwX9hus084BRZdo2i+DVgvXajMrpfFSndNN7nKxA2YO06tH0bvTHrTTkGFwQ
Pekyf0YGXJUJbg3FmS3d/iBGmabYttG/Lnj+eCliFE2AdauiLGEdh+y7Uhk8jHCF
CkeW7ANVL5QPnEWYu5gwx+YOFL7JGm/vOxk+QkbQfnmdixYVUmPWJro8L/F5lAiV
EkfvpP2AMM5cRpPdXOBJ1+aWyr7uiL6Xd7fI9EnlVnrFlCVWCA3X4Ut0piSjYBSM
sS2WOV1M+ExqcD/PPS1V6EvvIXwYn5vRZUYYtj+5Ju/xK1mBNWmwJxO3bzb1DU15
NGBmLu6qGZUKDrxNDIpzKm8yEyhyw/tGhICDya/DIzVJ7nz9jeCq+ZHjemj4p9ts
JY2TKAnZmh8OWhl6YvHTpn2JHok2dq6KoNseaTqelFLGxuoxI6/H3cCxYp5Khed/
YF5YrWbM96qW/Nv1IflpTzS1EEq9q9fL2yi8ErocG7Pn3jvcKTYNGLiIYSRcZSoY
/yxFnvGsomJuFsIbb7eJPOI5Hq4GaTsiK0DjEwbGORYVkdNMvUFzSV+XBJ9H762z
hI95Q/vSN29wAjeEOofp4YE3lse+nsO2RMI0llIy2N4lSUBhiYsWnFXNbkbl2o29
tKrk9XCHApVleKj/G3KovjRaDAJu4iM4DNA962BzZRe5FL8Aesb1NW4XlZIjuWce
BgR2xWOMmPmVFAVEZ4N+U0dujBS5UABZT5b7zL3076XRhdXoSeHKc63DLdU4YlG8
WdOvmGCXaAzicosgFo6ogyjqI6lO95aqwyX3g9XmBDUWdLmClS/HTGq6IBziQhMQ
GXMHfIK7wBSsjUEgIMykHR64LR7k1YbfYD3q4a4dDwyIG/LXCk8ylq6m5kkW4qe5
gA46iMs+5KouTgVJ37UqUT+YZy556B7U0r6BYOCYSUKIgyGw+Ewi8ut+Ul1ELMwg
wnCAc4hjWY9yTKyVza4la935MhwZmRAKO0OvVdFXj2+RghHna/2uxwlbqyChqjiS
xJpNPp3X+Afr8ngbaZKAhxyHKOlsB//zDOOVNId70VnM2FUMzHAsFliGsY3Tm1mS
FcIVrLPA5rE6b+gz4gGBYvukCFjsC6IcwFQBZxPOXBjNHubNrhnL2XI5iVIcbBeF
YJC5aZ+mmFlhnv7zJ2wb7R1zQSOI2a2HYhY+w6W/XqRfF0KAdq1U9bMv7I/GjSib
SulAe9hmYUwn2tF4Qwsx72PLB17qLgh9Z+fvbkG2RBAfS+/z9n3cH1bm8BPk7MQn
eKLsn38NNSEzzixHdD33ZYWlX7QV/HTbqnj62Rngd9xo+Xw3Su3yaSDuqDoXF8p+
WwINoGsTOUd5BcicghlM99YVjTo0fO0P5prBJNl3R/cjPSMoZKgcPsWeJlmV0GwH
dbnCgR3d440NwIInA16uG3l6RJnOHLjqzHtPjr2I0IgWWeNJR9JJc0q4y1ydk3tM
vC9UdIPsVz6jLjdTyuUmw8nuzoBCAY7+QBzTApet89biFx8v7txJ/XVsFQ6MxOOp
7UiWBWL9/klbIDYTdKyegAXiSXc/Zn8ktX3Wr2+r3GWwKa4UX4yl0mZwkVqOtVo3
nvTLmtxFmCfvctgqrGi2sKd2r5XsOg8p8HGCi8z4r3ALeFl6WrqzQz1QYF7V/F05
3flXDTGs3G+ao8iO9Ntcdeel7O5st97k/vnyW8oYEA3bLdlxVFCfgC8znznfqrpY
g9igix2ikGhgJZhL5S08QDErCOsAz+UhlizpgTuI/ahzICkS+L2dS8LQmi6KOFN0
HSuRaU6DqETtsx8m7WJnjkTAPTCTsiZeScTMZWP23jBf0AAnGZbxVHJ+5zS6o9FP
OFF3Tnx7k8EcfvQ0yVgGJVVBJxSPHJiuo2iQTOPWoDnZ7km8sGN7eOguTUXIRCR+
Hqm2qWL3H2TQm1PN4Oni4QoSFksE3ZT0QgoJKNKZ3xykEvXaAmWONa+oCsiYTzeA
KtfSaFD8gLsXnCtbfb6LJ/Vu0UY/suOsHeEiuwVbizRr0D8odjZtFK+kYj99AQra
ACm3ES6RhoAuH4KHN9wfigVaDtovfPFQKU79dOfZ/Sud00oRsTP6YvbXhkKTL6+M
12sWsN7TNQZosp/LpRluxSZTOJ2sF8iDKZqVYdsrPWzi3UeflLYpTrxs35AaqwXO
tN8kBkyTTv+HFJMUJxauKwJHI8q70lzUFFbLeJdqskQEj4OxhX2gADiC/NIagHPy
p6+uA3rh8H3A/tEpDhAABgzEoJDAr/HiA4dTjs/BibLfo222iUzGnra60uPSUO2P
FqkhCYVZajxlZcoCfMtmXLNteqMqZhoaWTEctKX00ns0WZVDBo5RI1ciYxyQrj1m
sxvHbgZkJNE2WZTGm9FNUi/Ca4aQSND76PPgxjZJkBtc1Pf3zms2Tit6DYJSN94F
kv1dJS9m6JnSwTQWvY3JydVjN1NmSl7Oagw8YfqqXMCndWhdtaNa0lkiDXwrEdUA
X3BAll+fG4kMlJ4ZXMilAT641VWKVo+cvoA5eqQoqqCIFt0Aytt7uI3iZ+Y/DvCd
mm0KF4bvO6wgNftyqLLp1RpEWvPj+LQEh2w+o89RADJZIsU23AdgpvPwYtkJKXQV
Gftqjo+XcS+H73sRYzhBvs2azcd43HRXoitmQpsxv+zYfw31WhwFVA+B+SO+kAj7
bZSFmdxLde0hKJ7UosmVNKmCd9z5XnlL/GVYv7lcRSI1h1WoIwGj6hWNB/b/FNOA
xprSldRCOnk5BJhv1VAujrY+U4J3LYVIYngSVyKTaPpNuiddAOwaylFxSukSsPOd
1BjHuon38idq2xTkWnm+yRMzRY1vGbNZFnm3cK1KgkbuO0jix+bPDigD4fwZXb6h
7GgvuWE5Y/12gbeFTx34Eq6DRjUpFpZieN9p299tKIJp+ry+Z48zIeP8T0PuZQEy
yOVthyaUnRPuiB2LZzXZOCBJQkWlsD+wru7vTeZ+/25UGCysLNrWPVjHo7PjR5uc
7gB8vRLly2AHLBxyHbhE9Wqf6E56QeiTXp4+StDmQayVhvCBQPWt8Xk7fFMMG/0Q
uUHWv6R0Kb8NWiRMGsSvEo1up6o9CFIFm23DGI9WtwXJ5A8ZhVBF+mqwb30sKw+0
1WlqjdaEnU/dvIgpaMhDG5OiwYRJSLP2zyePPGQmZrB21IQjs4KP2ev3doS3I1mq
kWw7t9P47ete9ZnIlJTrYISzuaywR/4sRsslUARaqUhxSjnZWPYP8JEmvzCC4KXd
ujjH/EEW6YdKKIW6J3JeJJogmR1K3op6xRN54Rfja9Z07OQbIIZ5HBhz4MbiieFN
yw6y7uoPT9b/NEDekUYzbg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
L3Ty98evxbruC4Fh1Kg30MYIeKxUQPwWg85+vQL4X2EbMbLbsj5+MfmvrGBaVZB9
XQmIXlK3VUinDNjABw6Kx2nvK28TZ+Rvt9HhYffSlwNT3ATDb98TCxmmZIZ8z8I/
IDhk6r9x07TblCXf0UMxwzzVVYQ1b83kdc+OvQ7oLQ2pKhXa4IczDu9mX8PM0qE8
k3SwcnXdDcZhrIGPOxhkbYFVkZVAlSZB/tkVCCw0SYrZGIFQygwGk21hTXSZ0olh
UaOrIRj4snN7E/mMZ/hN+s+cC8BKGRLjXYHQfWx4v5ZYJFDuIzTMxTjdxVM3QrXn
4f7VIJ09ys0g5Vakqbrdhg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7408 )
`pragma protect data_block
iYjCCZNmK73/5Xyyzl6I0n96jYecK4B+yrknkJMRQoPTbJ3xUGBDgczDRMW9TpNe
08FgWoPx1KLhAwNkm9pqltPmiCdV6UyqX6sPQwvbRZVVfr/CgP8qhGG53XnpeUO7
NcA7soX4lkmu+PMYevWHuq4gzwn9M7z8LHqHkeFDccXgVizt/YxSSiqkReYXiZZ3
84ilEtsx8/BPjU05OB5oZxArCHKwooEcRKlt8hCU4KtZJeakR5Lt2+2GUtZ64fab
TEB9fyqjH75RMSFd3j9pe6VeOYNF2BMcVSWXXericWIkwqzfvnkwT/yF9nBV0wLB
tKW+p3Awmz/SsO+2JCoe8UeXXlGz537TZ6qB5PDz/VTzXa4BdFoUIOMHhun+sC0p
63ybbPGVD82DJXoB7uAkMFAjCal9ERo5qiGfltdLyOJHgatkuoO9oVs/Ilr4KbKX
vehH7lVDtLUERW0zHFnFwR4rJZ/cbyVGoTTICZK8SjlF94296Ry4Qx/BMitzFbB/
ihH1lxRP9e/d+1j18Cdczv2UzIrYK2M1k/y0WqcVMknZrypsmUhEhXFhjt8efvxp
JRdvhYVmKEncwYbyrxUmyUTtlasvDwn/RcUUSejw3z4lwzFjggagYOoH8hnVIYAo
xQ2rBsW7TZyEO64qNxPKJJqjJCuVjn6QbjKduzVtRXglL3EAqHrMkym+4ITJIphg
mW8P3zvgY1SwRyXswEi3BzgSbVdcgpKJBa/VHbYOuSgns8IBsJCefmfUN6n1Yt2K
hbFOUj9r7egjIFfe0Ccoa23cjMWnVgSx86RPbcRrkZBTHrhJCU3ixw2xCKdvYGNo
zp6yzYYUR/PGIysufCpXyRBRfZ2XTfSu4/JJTIVHMaXqKkxLX5BmZnOTcTVTnObb
GHBy3AwZTNct4uJ6CUYr4HsbO4MZ6skQk7ryGgoZzS7UW6+RIuXXNMlH4AlmfaPa
BRMd4nFm59ttnLRZJ42+aTRZZaUvNmtmeyoWO2Nm5ylGDAeYErngQVnspf67rDt0
7h5k1QWqrVofOG18TTCXFhTFv93YW0U2MNxy6muRcOBkdsNEcch+Fe/1oVNb0pSO
IbdeoLPLl8BQQ4Aj0cWIflOCb5zM52MQD0yTo5j1dijl1idNWBDZx8IFWXUhcc+t
+Dd2qQ0OEjhRxs1Q0PBIn2iaERKayWFjGNFPdtg0KVf2oCZjedno6aychvx5tfBx
ftT0HqDBlSiYqOKa8alT5RM/hm7fLQOykI1R3+1KD2r1MeDmgzG+jcuy+j5zc7Xv
pAcqrsp766FUeeBpjkwFj1wxNdJGSUER+LDzHB/8anr4vTzYJSqu71yP05z2ME0t
fD7KuDoW/rxraG+A3nk+VCzVRYmiYViVJ+0N8dtmJ/LgvmoPb1dfcdEK+EmKFqPb
meLka1kSglBGUyYGKEH0ZaRnCJI9XuKyVcRApxXVgPPso0/fRPHJbEOBT6WhAxh0
gywo6rk3EGtB1ADqvPRjKXLWw+qbqVFJQl11nbaCkp5/oGNtJowGD54xtUgzFgKG
D8bD92xEmVMT5N0Hi1U1pXxFddL8racx28O+bGZ5jevp7WQa+gOknI6MzE94H3Et
E841+52NSBIO/oAzKP3aaAxHxbh8dh+nnxzds1uyZS1fBV9ai1xAiyqANkXTMMMI
lEFj+RelCCeDB65W+o1wiktZLp1lmbIJ4QgZhrCczgvybsn1SKl/cdmU7FkOtsRj
HLXyF5/RQeshPfDJaCpqq2s2vJ+oiwT+c3iBy2+8IVD8Lh2czupxRa+16bMEvDrM
eNykUyTvuyLVUljx+wl6bnEFNUVcb+HpBsnTMyEZAxUeIEe6Z1sY+NMpyolfe68k
KEBUQH35hgr/sz6hV+Q79d11v86BLM89aXiqHwp0mZOivEqhYxiyS6P/olX+ld1A
Wjpbv6kRmb/41YX1+xZ2YNNcuG8WGxuaQysv+E5NWD6zZOI0ypTWCdiyOsm6egXo
9GPSgP9l98SCohr4O9UT4v/j0sEhtm9mgg0PV9CqxDXM6c8H3cxVrwUwdqn7ef8Y
AE4/lTtKuDyMFDOEoqkcJVyAIej2tGJh76Qj6K43VWQPnIrPXnOL9ppfWeWv36MB
cgbZQspMEQSbu9qnqj86aPgHNiCs4XqLnKP5csLwVmVF0qSJGxz/T6u6EDy45tSQ
UUWrNwT3uTci1w8AJQSLd9M7MpskoKSjILlqnJZ/e4CjI703q6g85nf7flVLasXk
y6SyI96DYrX0Rcs6yYq/NCaBa8vdXkyoesdwftiYjm4j/IFclAkIowzYe6YCrlMz
roJYXHqaQB0HCQrIBzpKaDcLLF08A3d4I9GJMcxKrGOh3ildN9c7hH7IJ11npjuB
IZjHCDl8JYZwlFnAwFGujl72b0hbrWaPLiK/ylkZK0EyBKL+1dvFm92Ivzxw8Que
BJa9hK3QRIP35v7tNAiPVFXX346Bl1lFXQTGYleOnhB8IRbjaK/mGYgh3pF/KxX0
7rAx+laZ23t1MaSLB2ZQlkjWlVYLYbP+mndw1ylXgN0N2gMe8o6qPQ/nvL6H2xNt
dZFc8UxXBxf4VcfrGYGXbcSB/7EGdAGIEQ1lfMsiiRGQnMtXGmzBMX+AGIgQ0G0l
Dsbu9NFvwHWfKsU/42yZMmycH6xiIi0xcKTdIESk6qPqFWm6WPpqgzgphulEc2Im
7X+0OaScf5b4utqBfb/j3Mzbov6YnN/VGWn21nY7R7DjqI2zWgPkyoWegLDwGhwb
Cz4ngGchs0x41pOTZqrllqaKAsJQw5Pn95tEUYExEWXN86i03tVpoenDiYS/mmOP
TSPvt61RW2WFCVgj8rmKCK4mILXoBcgN6L6Iv2qgDjaaPyBsmvAiQHEElX6GukVC
W1C2tgst+qyxNR8/apHy9aSBOoR/qWEzVBx1/9BBZlYXa9OmFw95am26wDWpE5gW
FfEuwRYVvkN0kW/uv07/RoJV1nRoGyfcFbN42j+IiFtB0xhArvo/bSwy7lyQIS6N
FR4lFu0S9WW5xZ+dki1dHeVfm53kl31Kq6FTMyTbv3DcLgnll756g817KbwTKMCl
A5D5MEe/gy0l/lSy2OW3gZorVhPluZnhz2TVEPj0MtMpwVrDTNf5U0RFLLnSEKW7
3L2Os4oFcTxt5PiClRjPTV5MgoaDHqgEBB+JBGJ+Ijf99Sx+ewfk8+KxaIHNUz7j
NIWcCadkqgqVwyll0ey20rhA+cAmjQxgok8WCb3pnp2VTbRh/wV8iSTnlEkFRpvD
gO8nqtGqRCTxMl5SxIzxvNLfMrMPbo2dGZ1YCyCUIhPPzOtAJvyOu2gR77+c7Hwg
gix4a6nlsoOPkXI7ehWj/+IcNND5eGLXmaAFZTs111a4r5LL0g6PfnVif1822elM
1Aqcfaavu8/yTWfrB+LDvbQyE9IZQ3WYoQE8ZpeLzPFxiON/w524pi3Z/N0MWUcB
IgeYVNiJAB/B7mSqwmqS6B5IGQ9imBEuVDQEzYXjmBF1EoCM3VWUOcBz2Ymn0mXR
x3LRqO7K91Nrj/9XdNfqjLtr9JEnKIjYDvo9pIutjgbtRWbPEINyJlem1LSH6lG1
XUf3gn9Z89/Rn9Ob7G3Ap0Vm/qmXKAY9GoiJ2okEkvzukjA29RrmmECNnu5r4CXR
SxzJ8gnYwAKW07l5wEobGuj5lDcvqA9UHmxbsv02qBMASGWnVRO4JvliwNYUygsS
Bpj0jt+cAAsrc7ZXavj3h+6p0gfA1w5t5r2rMX9nkprRAr7Tj9mxYm2HaKv+qKor
h2Bn49MZL7thRHg3m3BfQjAdTiDTU5mqW7V4INX2qZ2tc3jBlPmKnPCc/Us+xxuK
IbvoOiPhh34iDzSpbQ2tmDD4xZcjhM1V15QBDyxgXRRh2R3b7GMHRjcj91ScFJ1t
/P4sNuNqKIkCihKYKCIX2et6MowuGYnsfNcoNuF1n5Af+t13W+8OlOLUG4mJltum
oDxoT2Bv5jUjJhUtUMn1zchu1DHjnHTo1iQsTON0g9Ka/GLgGDqpqWywxpyOkJLv
hcyUcn0r18IjaggdP/T1b1+Hbcqc76nWWaCIqHzftNOXWsgmrReJQHLB+KIE9gLt
Om5PtOmnthwP8WCtudyIB2iLgwPGVdGQ38y629qDIsr/ugZRclW9l3IAOHWixT0F
CC6LZbZM+2VBm05Ts80bdPuwgeA6jUj4gK+CVRrjqMmjkKf8EYV39bFi4fXJtbKl
jVCdUQMgTKIehLtgsL/nxVEx12qcsmasUeX4i7ui14bIzXJovZ/ETiR/J+OY1AV3
4oWwUBSr4QIl/d1GgFryu0UZAIgudJnnnQvXiykPTAGTMVzhUXixuxy5lOkWN5Kf
roAJq3JcecdP+RHK8/vlBolHXHYF7br8OK+f2WUdYyRhlTn/ZEb+N0O3SptbKyVQ
zPAa1njtpWNPrAE87Cd3mWYFE0RoQFuzcRK4U3OA4vuRQoEw2lOjO4LM7SFhzEfJ
nnTk30oRmwjvZZQP0AnsNMc2UTHktypNeY/XCNXzOKFvMLBkywubwuhakrx19uwB
jfRqEouQWVDf166peJmgwAGe61HXEhLB1llOUb5FNKomMeu8msRm1JJg40V25flF
zYQNCHQEufz5x5wO31JZmidmvHVDeP7gEuWixJ0eFnQDYMzJH0UC8DaSYV69dtnP
3AkfHExpQFCf1DwHY2gSCtIekUQxRhXkAE8W0yVXr93KZzL1ylbHsc8anxunWFQc
fLGH2agwqFnfUgM3jYGa9EnWsw2jAwdHDpQAefiSvHOZHDX7Rn5ZZPEz4gEI2ZIV
B1duLAaw6FCRyOez02Ww+06znbOMywbOJZsWeSOIu6AnCJ4a0+EZrtjJC/4YmykH
vl4H/To+RhksywqktCjNk9pIw0MbSS+Iz2TwAhDP8l0C3gnGYx29nOCD1k7URRT2
/lSxsUIeXLDR0QJgJmovQ9ZCUQW9NNsnvbv37/tWU86zlBm+RN2qRPT/MPpTrMzv
pDBtTAE6oaIvU2l0VuGb6JrY2qYRqPQQjEL+yi1TPkIR07Imn+R5t56OxpTtjccp
TK6d+UD+X/4oASOer9AQEariGern/V+utvJX/hTgN5dWR96zfr073rBhuIm3oIRK
4Y8dCuuDSRfoO+Heo/squxhh9inGmEi2hPqs+4Qp9M+JjIfDZs7pW+CjBl+yOpkX
X/G9a6F8Gr1+sfF8P0vW/G3D0L0Q5QlpHAe7IkZUF7AjO6C3gFuia2jNrPjNMZuh
qGeSXYoVO60TP2WpDAC1DyVVfB7jNSyyW1KSEpexOUJrvE3/m3QyiCv5J6XUw9iW
FqN7EcvZk5TBsN++ySazbJV07yGN+E7U5k5yqnvEoCT0vr0QRga5/l+1iySDjtrJ
mqXZzDyh+yGRsEEQWfOCgGAVmg5dP5JKHB3i9KhdqZIoqAUVG3iVbA9R37tb501+
efUT2kYqy2qMwi0NewnrfOJahAckn4MhZDshPSSD8DmgwYsKTQGoXiGRL7z4gN38
43rdGhe4DQ1iAmemJHmq+MTdxSLeDmwUyV6cWC082333SaC7SbjQfu3+7CsYRul3
PiwR37nigtA0iOHgt9a4z+totznzPMzEeBzejH6O/meNB34qldLNFACJ0vJhsRmm
A0a0lMTSHL+OhzC9rjYwt4PbKfLeajEC/UTkp6X0NL8e8TE64WdEi1z5xP1JLkZq
cgNGI1T1n+SpeNyDjUhTdMBcdZgJyCy52tqiHuuWXsbjO425eSdv/YuHEWZZHSrt
xH5SEl1+BHGkaGQWaS5ryx4QE33ZYuxSDM9JRfIq8n+03XJqeVHSiG+hRzsoSwaX
F3pSmW1bxy3LcvsMdbi6CETZQ8haehXB0xPdryVwnPuXyX1fj3EbMI5qIn0tgj2a
gZHcBq32bkRj3r2lvcDiJBfwwUdi4FZGx2Hp/VA1Z+LKiiGnkSqERf76/1orOGSX
EUn5GRlp5tb0QvKIZB2DfoilCu42WyJxCy6UoWG9ldhI8STTrfwYXTe1qXryZu0N
dAaAtuZ1WtXyPbiblUYkCST4fbtRe2Obw17wafdRxfuJ6Opa5Ipw0SBHrIcmTAmr
37mC8B8SwMu5Lf83A5q5tdGY6Gq96s56vSG5n7s230LKqnIH3PipxbspyA4zsz4W
lEdPnoBkY7v4L2Jwh/SuDoBtdryBf1j9bNfif71P40b228vzdzGi6r7gwVb0wAeD
3aEt6XcuOCRnUc0ezBu7qD/zKnh/pVK+2b/jodkhhS7VyfU8YscuXZVl/1nHd2+Z
ISzQ4rrdR44gm8hg5txVm3vSL5tVtfHcQwxnM0yXfWjOIAFeX2JcN8M6l6flT/xu
zFP4LqnPH4iIICbWDtdDjlOR8FPRIszkDXZSvRUvns8P/Islx486gfgTpiszHjBd
rayRM+IiNx/nEEndHR/dnRnlyBactEhB0J8kP5dCg1O2f2t3fA2cnNnul91IrUK8
vrlQmDbW2BRyUvtqNFFUyq6PcRIMUXb9Fj66pgpElXMbXj1HKFqiFbKeVklj1s2I
rV6Qs3j+4M2Dhk9RoexcevBTFuuGrKa2xAe3OMwglFJl5TH9OodHatlSivlXUpHJ
Ziwjecr2JqGE7yqGiiQtfaJIiR33b1YP+3c5wEdMSt5/zbjd8WA8D2zZNMba2AWb
oUbLGjIPT5ICVhNMVJ/9TXrdqvaYxYBCYSUfEaBYh60ZcfHi74vb5kPJQUJfh8W1
kn5fc94qF17PDhi+SgG9ol8ayvc7wRr5MKR4lEPXaUiSRPE2PNMQ3SuX80JA5HjS
Qcep7RpYthKKoy3LKb4UygzwOTnXvsWqXKz9I35vPUzoKcKuTuyTm+o54kYVCCJx
NLOECBpQ0f08eNIEqf36ve5BN+2Cjr1QX9BzVd/yNFcSn1xTT5XBzfkzDvNRHkV8
Hh91tM/I91mDL7RVMDQ7XSzVv0E7N+LkTvAq8fdnugrWfdb8jVL3Ulny8mib082d
chy7TieAD6B3k2ayASb3mqfJuZ6GCWstMaf5nEMkK+za96sA/TKk0EPHNe+0pok1
l6Y7R9z0I2wj40zqrjyUgEq09Z+MpI4CIPej5mNnCMwFQikWYh2M0EUrKDOuvomm
jNcDJ52OlzZaPRX7eggGbTXK0TznHvAYVTvBvK0oM7a7VyCju38bjSbOjDMw9FBK
qRFDw5uC0d7F+9jTuAefftw85JtdItE/QHr77LC0TgGYs5hXctolMc5PjynssRoH
jW88V/533JwSV6lJBu2+Nk//Q/4paNXXST7lGU9D7oxlOIYjnFzXUSSjqQ+xwMb/
MAyNWJzSoXarm0W2g5lN682MOcUBwNoJjH3SeepJtHtp1U8qwj8eRbuXszUjhQqV
lQNeHBPgjJcD1r21yDhsXFqyZmej5ghWjYFydAJc3z5mGyI3yLiv1/5SPBYsHPry
1r2qVEMkuztewWXVHWbzeKUijwblCXzDPy5oim6p0jIBVl2eoEIxxjOVF1Z+sKTn
7XK37FqdSyErAgTn0W30V2qV9+96v9avLVpke9tlbHguNm18rlsco+l3HK5QCXCh
408mCUaxyCG/bINowDLnOXJoM9Q0GT2ZZhxAPD3o+dCu7Ycn4K2P0nb5ynkFzUYJ
D2myniZF9u96C4hgVAm7CyY+cugeOJ1QrkT/TPRKF6eW0HqOdFLt8fKPGsmNocbQ
zlRzrjDMnF6Y8jRANQPJPVexco/6u55s7/XlpeUGMr2sDmNvfG7neMK+7YlmEkz/
04XuI7C+BtUTRAoS+Bb+TD8g8qIM0vIBknC/ItgjMXwHr6mcBDjstoTUSSZ+E8at
WQHSz0hMQzQEeb4k1FytfqFy8J8GO3u5CQua2mYJGHRL+UL+W7/mSUYHuIHoTul7
9odA5YmccilnRUQe1hH63T49gDnMcOjsgT7IgbWwlwCsuspD2hSOMS2FhI7YwWLQ
PoGKRGlKkSWNJr1pPopjxkqOzdN9kGsMekH8lmY9NjbP/jnpy9F7wi4lfgVYCgG4
wxf9sRdjZkbLwBV5ac8yfMUJI4/Cve1V5BP+GCd0lyCajjkv8upPg3zAZAPQTXUA
MXBLzaIAwT95/OX7ON76Z4kc6KUNXtsYPZmku1epPc0yzjtXEnDqoedDOpNzB8KG
PTL2c9XW1qpFpaq8+uCFZcrR1yKqKC1Hsmuekxk42iGQz0K+MrkhmE4/uzHMGfoB
pJyPzEHDlHSkOSfd3MJ+MTqsChX+CCdzakK5ppzPU2wAQ1I1/OASfcS5ez5UAmGV
1z6WTxouHdfwFELtekyW6mtGaxGL5eyKxtxZtUA85CnoLfTx6el9pl7Zavzfw+qP
Cl15sID2tC1Ar5MzROpg6euTcGwUJx22dAkp8GCP70JcvX1G/rW/cmCHHFMxWJoS
DyB6OTbNGmJ7mRR8VgYADRO1LshyNqCf+Fal3k04iVb0SRuiy/N9AOEam5tRvVQO
MAD2wSNGZdwQQrMd7TNU+RrGMg7tT1R7h7b1Hr6U4+M+xXcFp6mJBj/P3oKzUO8h
OXK3GZ2lR0mdbieGU3MiCApnxxJ7FvKxdobT3BrDd9UZ0DdusVHFce+9YVfs2Civ
Js3og3F8BxgXfPUd80L8iGMu27jA6hMm4y/GOSy222L29IHNG2kvnciUcksKv17o
M9D2VKGzP4Ok7apJezSh6U1XYO7z0QsN47zDBNoKFElNhuXIaebu2Wrapva3YDXB
40yT3LexOp4zjgBXvTmArmwBTBcDELqy9+O1oVFLOVsVTSDs0d0K2HnfnWEboSjz
YXd8Z1XfmKWGAHTXpimkfOsZScONqwIV1lKwO8v6+VP10entBKW67hgtl8KseCog
JIXkOrNcevcGN4Zjczy5vHMNFW1nIx0YEXg1ky4EcKPzvRqvSQEr7EfHf3JBGt7o
cFrDYmjgvFbHWCyUo/Hkyoxl73RMGYjQeCA/7n3njhAq23AAiOE2vNCuAR0bOvc0
SC6du1nuqiphnotvsnHU9AaD7kAuOAMdnjinNJ9d2wqiFl3bmMLjID2zGRtgxhaN
zqZD0kcrvlLDZhvRQ7TF/B3dBrCKS/8zpBYOy42CWq19i2saK2BuiCR2Rt7MdbFb
mAj7Ry9cYE3691AeLNT7Lfmc591sgTGyzkbNI0X1KUAqNczEKfP/URwVOsbkQuj+
3oBf1MNg0U14NZmUUNk6kCpzMrhV4rtDEv+7zUAY3iaV9SEJWb6GTOI1xuRkDJco
i+Zp4CplHPTAuSEvMv19COZdH0A0E6bV9YoTGGYEkLMKwIoY7BTDV6nsZRX/8tMX
ukcTsZUt1DHdEpayl7fsvACPD2mAkM2WiDXK/EYpF6cvDbvppQwOzoLaA/3an7fB
5DtNf3PQGbemben1wCw/oetw2MKK2uRSnyMcAyuH7+s2ux64Ttvoob2XJ1R2zsRU
UBTuTPgTdm9EM7a2ZmnOakR/ZjVDLPPM636n1g5mQ3mNSSJrRw0yLvCkkSr3lcXf
N9b2SC5jXgKEZOu/LAX+4BHvyRG1G5LBwF11GgmsM6yEFVCko1LldmsrB7GJHhSm
ke+9Bk2AE8+OSCEATKT3FUt8uosIMT5zo5kdsmCL0z6ohzV2HUXzEy3lqhpLTNfb
Uj6M2z4OC0T08D1t92x6vpL1y2181JWwayTVBezZFhT+oXF67QVmTF2Vs0yD5XdY
sbBAevTGP/V5PWUlnOBGcmrYlBkacklEo/AGc4qDF50yQou10wl2u5ebjjyUTPNO
RXOH1DL1viKg/HLtgHiEGe0DLcWogOW4uhWojvGZHn54L/J3yWNAVwyWdSWs5VJ8
2eC5JjPzQRrn4jPiFetLeD06H754NqgRPI1R9wkySfSc6pP5k4J4Wx+e6/rQ3ZJO
cT1AZmjqZnlO2TiU7At6TA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
e8GX9cDeV9oBCbz67nDcgNrdvcxMlPrJDiy6xkec8EDaQU4uLyKmW3k7DFpTUyR/
+1+uSKxURnJu1FUq5nWzJBzJ0pjRB7vUtgkDVObxN64RYZBZxKMcxJDvinplS01a
wCIffM0KhNELAz99cIDT+YNBzyYXY/I0jltWg9pWpSKqG3TmEVB4I6310y3ZjB9k
Xs17oXKGiMI9KfgWIV8xOBlIzO7BIV3yYFRzddUMh/VoYkRm52glwFGmILdb/1L5
2+nO3VdOLvlLzb+DX1+a9pWpyJYVwsSfA+U25Kiuhaiuy77U8fJvnZJeKCzfHaxd
ElROdo+KkC/3DAsnLA99Iw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15952 )
`pragma protect data_block
cRVLOb5OZq8wIULSHZL9sVnytrCz8Y2x6HCM3VMLnXzBQVEiikyabMTI3TRmkWOV
M1rp0dvNRRZc6V4H9WRvBOLj1hi8oYkRRt1GgkxiToV/gAXWGMONBUHQWypOQt7D
o75CtycUvKGFHpxuRGkToCkHeJ1RrLIfANEc3/WtPQEdjaAT09i92bXelRZqKSUY
xK+QNjdByEtxA5nkmv6HtLi0extyP0d5xZQeFGcHjvreZ2NETs7fZOgDtg4N8w37
eezc8hGZztwSqcq64inhaVN3t0thIaQRLLIOcAxZxYwK7haTSc8X70EMp14MBsmQ
ZDDRrdP2UxEHzNKRyf93/8uAE/uusvrjwElr+ivUikY1M9+KffWNOpyAW1mUXWBe
8oj3qsui2Tia2AFgrc4+7QSm16EyM1bIvelJptSb2xYMLZ7RD7FPTVRz9n5Fb1eL
WuJZFe2DqKnbww1hNoNxabrZFZS3KITG10hHvlpXse81LdfPndd7gGKQ+DbVKux2
46j/RWiABXR5CzNPwMf26/kRfX1Cv6AcTq0PCBaJOS8cEMqwzygtZEpQUl2PYCXm
l9ftDHayAVZlpsvpiNhtrlggxV2x2b6dT6EHszpO+Uremdw/vj9+7YVYTHdpft+b
zvfh8Sb5Q/uWYBFiIy4zs77DROahE8pJsHmicpwXUKAK7WGdjsntWy7FgP7c014V
qVZEchAMAOjlRE4qaTDUp+3jSieZbS+6pV42BGHCJcGk5XQH6wbo8lUdstho0QMd
orHPYwS4Fi7yISNPmgzhpf4qu54J6mlmXaB/13QBJRJCrXP2NN9B4DWsxfqRaPDA
TNoJVxzbiSXwH7abwRRIMd3ZQyBhT9yq5c7Yk0AldYJBlQUsZ66WHQPN+vjGnFUu
4sm81qQ66YQMyThlY6J1e83nxBID7kchZL1HxUFy6GCNMisl9c6m2xlmWRiqTT4m
ugo8OG2FH3F9jCMQGMr/nwwz/Q4EgfZ5Pav4boFbLZVWgTP+zWCeaUEv0g/9Msqu
K/IbUBmOpjYhT2GEsDedJLnpPm5emxtQGkFDb5BZYJQslAFjeF/WuVyBvbMh6kZA
iZnIX+t9/Rfl3+Yaakf+OnbBOxReAFSHYXzTMnd53KQBtnvSwJiHQMFwtaIoE1FD
D1B5yMJXl4wTCZ0Bl1zizHxWqtGgtCQoAX820TcwSEoutSBES6FT5dqlo8/Tkp2W
pT2MyejSQBQo4CKyZiq2yvAdTBmmA6kMj6AhJfMeUHqbo9VY1K4VbHcurIKrU25B
0DG4d2ftgvr38fjL256caWt5IaPvZufi6bkdebwPwmOERPEjXSB9tIcwAyPSNzHT
wUe/vjWSIB8EvhUVTneab1xuvgk+j0HMiU2fUlHKj8YmKWxCfLk+x+UICdcvd7YC
ZcRxekVWTBrYTwELZjSEsp9lN2nESap3L936RLQjiofMZaRbYo7PF7qdg2CBAUyh
poF7UhIntTQIRWlSO3S56vXV/2uw5RhqfjtCFSSNsWDOvmZJ/X1K739qp3EbKGPE
mXslmESGQwNDu3EfKSwGp2KV4apNbk4BVdqvVEJ/OTaaN4wSEi8ngzyM6W/7RqO7
bMYRR+rcgw+rhYuh5uEZRMFXAC9vu3eRRe9zl9lDwPcWsoaazUI6a0zAcEMokY0O
rRjdRDIvXN1Rwh63gwdONKd4YnrmeHqT1Py5FK4YG9OQrei1E8GBkpU+QyZJCqJu
z3JAacnP1BcR4iejxFQV8CfOOXYsPgluXtPRulEoqNwh8Y+zAEIEk8ngkfP0HtoA
1CWF/EhEJjvkf4ykvfJocubW4KY7g6DBnLFDobRaKZcLxiGg8E0mGJoBpQBpYw/G
nFOY6dTSpu82GauQs1p84EWx8msy4oSdhqPNzk62Q711/YbUJfTWROcIUAg6xET/
b5Sw5Jw4xRp0nkVmlHt6IQ4/X8X/6Huu3Fa8ELAom67LDVV3uO+K3SQSUsSK3jEV
jDemNMClsHtAp5dHDHH7bDDZDTmJxB564l2aZho1qldMwaSRi1FvsuLGsf/AI3iK
r8xW6SzahVnOq78dw+hTs5FdqigZN0TV/5Hh0X5uJ8nZTc8jQ6lFzNVmvz5rlimC
7mjv96wbJts1VHFdV7Rz98rLPhy8ZTNTolQc9hyiA4RoBggPijsXMhNRotczeYC7
wqSsH2ruggClduP/Ujg32lKxh9WAarRI6bZbv3sD/DZJcq2cj0XY++gGNMKoljgJ
1norgULghrxMt5FCW70HCf1mzYa9QrhnCsH76aXDkkah0KhPqF1zKEun2iklHytJ
VU0zAyYxa8HBrUsbWKLYyaV3wx6Us41YWbZ7l4lE6rOU05Ovt2c/bKpQP6YAV5yB
MU0C06OWCz4vQQVLxaqCn++gOxk8947wXwvRG/SqExJ/VPiOyjYVraB1ctiXo3w/
WTaKMptFigRW6vC5QGND8GiQbNP/e2G8Z10kqr//QQHAeCkxW5aN8lso7zD5ckc8
15OfClqifY1BU/bwZrizYYWtvPrdnaRBL83pn+ce8KYkpL2k6nblmZ10kFR9URH+
+VlUghpbvfvmvhyZGsA6wXt1kYrhT5zxIEWd8ZlSW0IAknE0uvO9V5PTD99SywJq
BqygBrjRHk0WuMKM+vRLnY46lcUN9aeJenX0YCkYm04O+UcH/elD1V5oN9BEjeZ4
GuSkv6xSz7P7rFQU+Sjnre3GBZvlD2pOBrOcpYGSQvpYmYw3soShCfJSseHBuWlO
B96vRSBaeZzTMp5N+sUyjBpnq4Xj+B2C8LjS0BuRo+YotMiTKT1+hOEaC/i2Y7y0
xx9zglgtTHvlQkNas3c/2OzgrAknIyuuVdpqUX/blxrjQPmEHifxbvdQmB2U27BU
O6CBHEH3Z0Fw5qkFYdf/b+oLQ/U3UgcYdUpw1WNJwF0TxYm9FIINjVaaWb7uuyQJ
pdwScU7/NWjle+bDmwgxjLwUt2hg20eWoxK1SxW+1I+ePIv548Is/n5wK2WUQr+k
DBDYVxuz6c1FkrReusok/kwOHT8P7qSyK7QmsgpzIStcORhxnvNiqIX6ZkdddyaT
PW2EvvVBHRktaZuXSe1IYqTGLBZoX5BhqAhEVev9A5M5rd07jRVaFBtiSEwTt66+
0HgjfzeMc+0NQsaa3wmxfShaKFdz71LAvrz8vS8KPH2aOFy/lHkedoHhgzzOohQz
umvuNt3DmUmeoFUrydjcfyqthpArPH8aUalL4ONInpBDh3pdNwWiXgCusHOhDLeX
eeUqYD69BGv65DnAlEMpaGRGPPbAN4Tm9GTdA0WnlqiSZgx+E/FCg6kAHpW480Xs
voyACvJSLtdBES6TrdW9KWr0tmSVChvA4rBZwAq2bNCNY/dLcoGuXefzhiG81M1L
6s0kD3c/l5TRXSlMrcauv5ELFBteA8SLO3NMjatn8l5pLU0NCooCTealezpp1Yu5
apO+IReNGFNnJrlJByA8ZTyK/w91d0AEVlZrJMqTyUENW7ZmkqoWEVgIoQhMir0W
ALYmJVULA91Cr3qK0Jd2iJPTOAHY9Z817UghRtn7/X9MxHhJqLg30HGlJ1j5fknW
4GCiz+hQjPP1I/JjFtBndjGSjDkrMcHUxkk8Wx4VVLqzmT01zvLO83uaZuqVn3Sq
KJFiQwuryBARhgsixRzU024cL+FgCO9DI80dbLqlnJeyUtbl/b9mqlDt+wGz6p8X
TnnE3Jx6feiS4Y9Nnl24AHteC4sfLxX56F1No80Iciqc5XhvX7Vbp62dX07DYaGg
52DiHE36J8XJ7A7AbeQ6NBkdLvZmOPpGVI6dojOdIvi57ReCWY5CsE94r3zYSfu5
eR8HNm1CKUGQtbVa99iZJkJGa4uz3VVak+8ZYE3nvOJOp0SVHIleU/kLpr4/7Qj6
+Kl50Sr1yNh0yGkaLYBBaG5FDcPmnY2WHrvhyL/5uanPVV95bP0IB+60u/OXBXNQ
LlWUGj6iazUfR9rmaV2TzpbLipkdrsIlTZkzt6kMHwZh/k3WKgYmJoYgESwDUAkR
ihyFzup9WCfFfX1Bf99NiRa/VX26FqkJC1Ua5K2g3zeLnXlNQtkUF3GnP7xvTWIx
hOP/+8H3NRykbcht8a/SV/gwKtTJx6krJSJwewVsaEcemuN+NW6nsDnWWbq1KgKi
6O8Ptxbf8WiiCYUSQ4a8PaQ52VrdCxmvvQykUKGpoKH1by9ntNuzXDvFi5LxN07g
S3RxlWb2WGJOhWJP+LIvKoizIwt4P1aSDtGx/H/gHdT0iMUVGcz1JN2wEYNeSUwH
mmYs7rAU40YrJbgBEMLobsHQnRUaRxcWlIi/73c/AlPReEUwXiNCflIPa7nt8Rik
2954VPVJ/8yAukGUsVsC6NHqZB0BEsoS6/8NpPR1tbkamnt9xvKt73uO9kS5vpVX
4BW/r3NNHRzUYaiCorxJWEe+9QM1UIB8XGduB+w93xQ6/j0QeuHF0fSZDyCuNnpV
YP9m4JABA1SaBOhLmtI9UfAAJsroOFdT1PDHB5bZKcQj+EPezkC+TSkAXhF/ck3y
GU5elBkpEp4v1143SSzWB3ZLa642mEQiwOJID8oADCbYUu/A4X2qFlpbHWRikapn
v2eay3BHWUQ/Sy0uA7VXqMzblwqPTugvDzyuPQzAlS5cnPhAVH96Z/DIuJw2ylTK
GZgSMDi2TI3vYI3x1Xkakk/bZ9jFwCBnwMR2gRU3xk5Glav0Otr4Xj8UF6sKR3Oa
q0kEo/rJGMdiuyHXibfzIxB1OkMEAZ+aOkp2f4hM9nj0HvSuD2hwkVWYpffjhbfm
eGZAQfMXA4Pedwoq2ukxCXyKubZXl6SzbYEBXDahDXPJS0JcE6POAsCTaftwIVyf
DT9GOoxWjByBEUn1kGfDLZPXu+DKw8sN1DVLvPnmttNh2q6yfLOK4B46MskCO/hI
XFx//tRb0kzqV6huk7StPkH8sdJCFHeZY/ACVKbgGfE+eekVd1qvQkOPveLBtBTM
lbF8p6fzOa4NR6jwqYOa2EGUVyj6PgMrbSFR3ZMILD2mnbe4oYJsxhF3RjH1wAJY
2dA2kPdtijoirueUTJqsUMweKUlXamr/ZMCjOheTyxaHpCFliZn2OB99hr2aKUjn
+A2KqOXU6EbQeKuMWVClevpv/KIMmItd1eydEKJIcQT1xR/8FClhL3jqkPeE1Kyd
c/aEBgMU/TGyxYEXACuPcLh6h6zaAvfjnmRKaAmb2JD7+mrLMLig67l8OWsA39qA
7nJZ4Pi/jkHDGQ5lKMwYyPCUPUQGKqNu+YZI0fLqNGqvT+f27+1ToXavHy4yxE2O
NOpo78snSFOLqjjjMwGY3sL631ZXMHX46G88HMyeRvAPslU8uwYYGiq+pS+0k6oS
5X17li/cXDnc0kDZCqHcFBZ2DJCUHxZUFZVpwVNCWZEjcgLvylM13f2jMe4V+1Nw
2wLQPkIV+kiSN5vcwgQtTpsvq+4AbSN4ftIBOE2f/v7S0o+ZHmpEJ7S9GOQoHDEY
tihGqO+A16vnfgttdTZEL9B1cEkTJcirO6mkcqLKftAutPu9R3hsM1kDbI3CgjEF
vouZzDiU7C4K6maGl/12Ci/rbNuyI4ip847PgJb0CDbfbMuyapIcMbz8le6Xpn0x
VUaRiXR4UNFc9ov9wsYiHrpuqkFsmxZLdLyj+0dDvOriqA55+qpd7VbBIwcAIu3R
XBNOZVAEVV36VlUMtDO9cgddjBWcPt2KizxhsbHQmA2EYHeJz5//M1zRCxcHNp+l
uvM67qc64MkJ3k6Lx3CQ4nFcA3vk5zTgDsNvgyqUCluTP95BIwpf8YCgyVEOGob8
FcYtwT3fl4VXjeKVj64zakU/j5xiJ3W2EoHKbGuC7rJU8ghMxFMJAJycXWfwdGHc
gX9D3l7HWvWcBkbQt0sFnz+BP133tGXjZbkMknmRyYeugzMh9mLpqMvXrCcV6rpO
SI464MRjjMQzkgfM0sREnUSD+NYBaG7O+m1+Ejo4h18GdnPyC29zIIQNQIOKAaIL
dWUNoBExDQA8oyP4n47SgWlMBnxqw35wV8V/JcoQeqE/mm3kejIRm7bpQnSVc2w7
tL6fIEnm+IQpuLs+I/E5F+cYmF6cEcAIw4txeGnHvc50E81okNW/jf2C/4VpgN1v
oviNp3YRyFAIK7n0O3wdCgcA1Fhibmk+FEmD7B+29Qf8So3sWhDqHn246eq7TQgI
aezj8qbSjugQSBEX/rudTDKxL8KlCgOTX5UdUSAzmKP2BcqkA42e06IlINJamcsS
UY1HjDFSpwjINvY76g+UTohz5hL8PrE6hptooHztgrfLGT2zfea3nSkZUqdEolmI
dmNO2wRF5FLqRT0wFIAwZftmQ9yxFgy2fo2oFYKvtT5dlcESUIl9qAxPe87JUDAj
bmZGvJht/LkW/VwT4awntlcXksSmPgmvXClo2UCPODQdRIyI0DV4kDgru6XBQhk0
C5puExOH5G0bWMsIOIWMtSjw7YwtqwwULYAE3XfJoMLGtYaTAacCAerdI+kfBQdB
O0n6ZvCQXWEvvmb9LXCZitSSR8k+DE7xIFKu1KcIbUoyyYwMaHFgPohwrX4sIXPK
l2RuQzTDfa+QMdXU2TJoYLOdxDEXg9fWY+ZoeuhxrKDWevf//F1Z2Cgo/CjMmq0K
9YmwawpxdfhL9XJYUhksMdLdtwJDEXXrDeJ+i9+wihodBrnGtup3BpbM1NUBrr+I
6eESxKCJPW5taJchfljjWhT18mV4OF8kr3y6RSKBi12NNqbjc6TImvlRjKaMcf8H
mdLnBCdznEGeujr5InQYVTVesNe+oaHh1VrL5JeNBjVX29PfS2dIEARbm+rhtxwJ
GwsHJE6Q84w+SUb1FC7AXK3/sDyZwVZrrEwIW1Z5ykfF52/uZmKGWkdCA+Pna/Gt
GRe1S8KXwU71RpPwy48ate8PltAZRxaNAHqtEucDhTO6fsDt8CfHCUotMLwJCgQu
RZpTLJ4rIfHeznp1as6ccgGMhltm87uJRt9BSO0AbNXxbbKhrRM0tbJIFpF5NXmA
iz2UDYt7GOHdGluVpGxAoKOPuxLBz3QamQiXD2AMzTcjHC9fox0XxyIK7EcA4oUZ
Oh+Jzvr6JXhrKtqXckju/m+EqUGdwlNrJrQsYfWgTnTRoB51iuiRkGBQTf4Wmz3M
Js/JWcGH3WFwsuE0r8Xw7lNdX62TClITgUzV+oRATEr5SHefyZm6+YeLQsIpr0hA
De3XbteafXsQOOhseR1Cv80YrBlJkpCxK3D6v1NqY52KS/t52Cl3uKPh8QQ4SbLX
0ROKPsa89kFFu5AfPdiCX6zBUGunIPFrCJayVOi0vKI6K111CqWpUvmqR3Onx9w8
SSUcsPheexzaD0D1OfA0TmnEBVUvaSToTSDf1Atwcwh7ZopVNFde1m+gv2jIn9pb
K2hOpv2+9bozv8BLP0QpxFQ0768c5Dr4qXb0P37cLAwdDFoOCJIbk9+zTkG8TFCC
X8geNHe6EjQCXrcrC//8xkfumGjlA3MNJR6qNG7cfxkW/4Yui/32Zk6WcVt92VS0
8OqgHGlan3HOwkldZJiLTLqs8/i7I9P0j3lxpN4n7Cag4tQJR5B+7j+BKqqcvGvO
o86ey2zGQbukFituGng7ah+Bjf5LQo1H7FDDi1+MEI7fvK4FuqCvlvzq0pE38oZL
pzGVhFRfNmy/aVK1wCT+dW2XUOZZTd0bC+7WBbtFDHiWW+J33PkLWAgPceSJndHz
F36/Xlc4610QSJLh9WF2Uto6z9yJkGLNbPMf0U6nVQwcOeRITk1g7XN6wWrbDwlb
4phswsgPl73TCA/O3MmDG78NpPCh+kGvXiEERMr/L9YpE5ATxx/Cvo5Xy5upUiXM
FEZu+ryjdnNkbD0lThlR7dJ465fj5pU4OuYrBb0CoZKyXOcbDCglFE7vtXHSgTz6
eFzqgYsdPZo3eotttSuC3FZrUj0hQM48mqSzQHTTwAtcCSQaiRWWmbnXE4TUd76Y
MI7oOaMIlNs3+J8Xm78FJdtNEL5xWi96GPmeT5K/tYRY/d0uFWexIMcb4b/gnIeC
jT+lirWsTz6SyufFMgQqG2zBfop4oRHI6ndMg8mbw3y/snlMK3D1FjN7cQkyiymZ
Bp2m4gPKj7rajsQgQN2eqzcbPxPwMoalA+5jdwDEHFQx6kbvrrR8ZZdB1xczWraS
/cFUSwNev4xiLzis2nnRmqPCQ0w0C9yPkzIjyqxcr3hcmX2flkWmvnwDibXzINCe
x84bWnIYDCjbHxKNAviNsQ74xYRs68BakEyVcNYU0DFOoJ6RRCFiYIRHF2C9UAFb
xFHHSRokCDVD+5amFU2ouU640T/WbrVUeMYuOrd1p1cTa/b764JrQAFa6nTlAXYd
gWZ3KSPAUgtmxtYPpFXffTmisxYbYbN8XbRIu8/LGxampe8vELThnzxOUm14O48O
W9R07llDpNm6EPFSiCk7zOPdR/IFI3LOU2d0R57o55Sj0IiSVikt34g/NG00QiOj
QLmcp7iGrPDum6ajNKdPP3OxhlOesZSaBDLdszcMsSd78wXnzreWtDx84QTvK88F
AXSRTsXW/6v0IpTsZksDGdJju7sOfKIEVKi5E7KKnX6wnyTSEcBTf4aquNuvg/r/
oMVfRA0nB2HwCBx+9Go0GeXNrdDiB6A+X8uzoqsgYFhXjo79Ye/x74ZvorwEU8j2
Q3OcPOOO+2pSMqYQMOyl4wPmZA1QulChTLvgn41XJQobaPMLskUtwpk2xUdzhU6l
7+0eyyZQsf78bUbUia0WQ6tgFhBe7YTfO5WQPpXVlFuo2tnX/zchbJl6Ol5lgWY5
H0E8qYgH+ffJILraqILLPpME3b6GzYlld+Ju1hIVcRH2jb8zngjODSsOqt58LNp9
kGIKngVM5SGQ9cpUFA+anWEEkeLOZr8J70SdfrS71X/k9e8f4i01bUkT4fZwTOba
VB153q+PuSkIh/sOGIGNoV9xDc1tbw/dDBRUn0CwZQFq/6PYBBaMNwswaqxoPV/m
g8Elx/9wxn60iUdGU+McgEN8bT+qqVmpnF/BDWR42VBMrywW9qfJ5KA3tax/835O
je3Tp4GatlgRJ2HjMuSUcjKk3pAUDOtR2jwMUnoTf947HaaINKucM1Ds9x66b+/y
ptFoHwS0Ydm0NflLgPsgF/MzAtauq50vsfn43UH2yXljPhq8rSJnZWCTzoy7mCF1
D807J4tIttrWL1tGNhhf7w5zWwSiOrVfkfielTsxaNoQ2JeF6KKnC4H+jX3DU+70
I0Gk1Vy+TUxSuUWpbxRVvb8CTFgA5DVedESef8w/anBmrlukChNiHv92aaTMyj6m
IsBRYH64myqXeub4Lzg6VTCQbBzNDNHGqEyYNMqDiKKP99527AU8c4UFaF2n6RBY
FgFIAzCYCee9LdAZgezONr+CsAB6xnYFOiXucKchUZEYspHWK1x21pnkCqwOGAzR
z/UVI9e0LpTZ2lJNvWcGWbBmXUe9IUbqkWAApLK/JsnC2G3QXWwHyWFrQOjZeZQO
qaheX5UaIxrrN/BIVwfWeZ7EduG2NOHPyh8rdTAG4LjSQPD6ZA1E0JhEfVinMzaK
ylh1+LbXRz9BTccQTZwGDK5xXoQo9qnX4BbR1eX7e4RSdxjTPl0jkozBZQYALR0i
GRnRsGfVeRRpyEgX5O9ALttbjU1vYxkBEBconkUbN7mYxvStKC5+/OakofSLxZB2
pntITjG+VYFH0oTeh5I2qDGGDmB3pWFeUe5X6kdgsz5AM73p2S5YEup9e3P2rvNN
E/o0o8Sq/R2h8RmtSEtPmdUq3CYA/12/e/FfZsZj075lPgZhZInO8/tX6uGc4Qbg
1+0Ry6hoC4DNwliqznl8s7MJdUNs5sMFioJLAmd6JzYJpD/UZ9GHuUxdx15Vmywt
YLXplHou+v1Dw3KpB1KQ48h9U6Q0H/j5Dk5+TrqIxk19q6HBpDmVvOF+C2Pe1EqG
KEPWNAKGG0iuRllimsqnII55lwLDQErlJiRccd1054kdjO6vjXlAC/MEhgGGA9nb
MWixpPNtCXG1QiDdAHuyakhuZJmrkjiq42hlnMGYnrhq5NHfgHBlsCMGzdaw3Elk
rODRoQjtWNvV/yh2BbDMacBCYTo61oKkOh0w0+LATkqrQgz7x68H0xYtJKxLcwOI
4ykz45c2yKc+yuCIkgKYFqzW46d0OX2RV8UcxaI1JM0kR3wrDkUKqV/twtlvwKbE
lrbVShuVqk50sPFI9NyRMZBeUjzne20tWhBOY9JrbXt2Txp39WtOf8TXmeXgHeIh
FQ65olcq4UKHrXsK7snION5pzzEmtCEp0d3OvuvwLrQL0PcWPaXwYMdwr3IcTNdE
NMYu0ZTXsZWtxmOUL/cQKqA94Tvvb7V1AL/aqDKiUKfwIfPeYZz/O9Zfv7LgPoUt
F8HG5Y/ivSn9ys/QcZ1zujn5eKszKklLjUQsdxpRHedKWIS3+1B0+YLV7hKPb4FR
NqBBGYjagKAaHKcFoJuLn7U+6+RLGModtoO3V6IjIzDSxivxU5WJWnQHF61DMCgd
fGGtaaZALcLYeWs2hLWr7qRspJQpi8CG3v1ph+6DTyCyoW6zPc1Rq51Zx8RJpmGU
hx5CyeJ4PJT7R/9Y84SkR1eZ94B5HOIteq6WqbJBIQ7CytpVavhbj8XjSh6ywLZG
XrfyVd9/2EJNqjtY3Zad/+ZFwKOzPht0Bl8+o06n55KxQykP5R6u1Q8tUfMJjEEV
f/nW6etmET+L4JkB+GVhaRklEzTapYZa6WZqjg12vMmBiG2aYykR25hPdHBsoYcz
krchqKZVoj9nHM7tluxgHvvMxB0QF3OWmYaDHI6HQ7aAN6wsM2Bu/I8Asax8Kdui
inIc+2IRlxupJONAEzqqa9EE+arlxTt35MBJClVHvveLxQL0kNw6L9oQ1xZ6HOuf
nZ0RYbm30htqTx0gBr7VEHOo5ZjiMxabK61mmKpvXqqa8yOwDvibX5TtjRjjXCGp
uXtD2M7//4Ygfgy40SfkRUbQnxLfeMzgymZfxGssq854vtGXbhqYwJYg2z5DU6uk
KkPAGrHMKycdzyo58nDQ8bv43rKJtKWZRYcbt09W2ilRcTHGLqkZmjfu3s87st9v
DxsIIPn0ClMaPv5gu5kXKbTXzPWmEhHWtYBTSPRq0YGFooi4ua+sDkxiQSovJXaQ
FixZZ8XYqvpPMdXflbw1dbGDRgU31G6TfTIJqE0ePAKte6rPUzoJeHaURN+6Lv0/
0hvxtCvjLHzexVaF8pvXMpEL6Awrp4LL34ew69w+wdEYIqMKWEjLAXdgwck+OHZy
DOloqC4QnMPM9ziD75sv/cT36kYxHz2CejVlJsoDnzLUVOn1kwSrLBgnnks81gLp
GQUd+UHrrYKUzPIQtqzye//gH0tHuCYdfCdfwiXnpm33iBdm6BGv1skE42uJpP+a
kW5TU1k3UDh1p/0TRGgtxeFDNfW7ics3+zE4qbhK6Ho+jjfdLH/n4Tg8BJgwRGwL
0fMRemDoa56MKUSYO0JlJNtYP+Dz8hEczMtyTwe6wb0k4WmGSqWLVhgQeVwOH+9g
sHP3l2OMqv4YLcIifpisnDlfLMCFISjzUsOTcWDIoaudP7BXW+ecJoS8SuXivl5d
5uSbLDHPpSl6rSps9Nzm8uJztoPBfTaME23Airf9Rr0sSAl1ESHImWCYgxi/hGk+
y8ITHFSBKCaM93H0Z09eWJzAHsW7dwpFStho6sH4e15eP+TehLKsTdG+XKmlabjc
3vFLRJsTLWpEMb5/DOgZWqwKHIfkEe+c3XoGzS70Z+4uluBKXr3uWaEtpney1Q+9
7uoeNNbqA6ayb97G7tePVOqKhyo2JWfigvhka9PZj/rAOejZvf39B//lO+QkFfWE
00HV3pLwqWWfd4+pD0WM2wzBVKF8z55XERxA6yUwDSUj4ymSZv+EYZyECjvqaCMH
+qrSu8QoU9UIlTb3fDI31AsKAoV1fy9bEJXhNzAT3m6d8MxoRmEe+Wlu9g5AQXRC
WaQMJfJxZPSQlml9/hDZ03r4JeZveYLu+hon4U5D1VLRUK302Kr1nuS4Nf5ueTGM
fVrOQymIIyaq5N4ypjwvnvn44IxB4PW1UFAlLB7ngPBE6RXvKZpexlMu6/nmoDmT
UDVhYuTr2k0vYmDeC0MuzZGJSh5KqnnXFHANCQDfzdrSYUvtuZkBjhULwsGIoZ9N
F/ip56DvRg9sZdC/0dfqjczXxvEXZLyqJKADjLyllTahy12qUpQB6NnJz6Z17kkr
IWkiZIdnt/POOserdxnSvtiu0SZrzvF5W01CWDPB0WaejWvxpVsgqtddqb99HIP2
2T1yyDf0uX+zCJA6Iou89uqiLJv4Qv1KFEe6s4X0RJYDcr0yqhkETeXxNzmtGvoY
g61JR/SBw6VMdC8ldCLILPfNQurQcuOW66pr9nj4jz5LrNkBFi3WuecWR4HR4/Z4
i+90ukC7IQIZn6MIWMNRNxN+0oa1KDtYw/r3+wkE9m7ywDGydpEM9u1ZKLdQkkZ7
MMsYUyL+fZzNtN7FW3bgeix0ovJVIntvU7pfYCENZhYCWYAuIH1sgPM6F+YtWl4Q
AS/HpG8EIA8RcFcR/pCOEeaY39fmHTqubXP/hp2EJ++chYqJ9acTHILKrWz7O8bm
T9HC6WA8dDbolLw6KUR1vgD5HoIwlHBPfuw7HOLq8OWdPT8OIKaSP+UdjbYONjM4
rXT0Olo3xkQ6h0gRgZofoCGINakK8wkNEPTvV8zOnjI4YsTykqR7g/UrK7w5g5iy
HFhJhKWOckBVXrHQxLUn44vx0yo7bpH9U6PFPXeRNIXv1IkigxA8wPODQ/jU+qmQ
LtzEgMq4JXUjIB6KiWb7Cx1vC/zG3+lk6gA91o+wxkbegFDQ4cNEG77VGP/a3L3Y
WDoawLbRc2ihuegmNDvDf9i7z4GgMxtf+kXoEa0sIBbIn0+AsyuhDSWMxYFlJ2Kq
mJJ0hOG/MO/HkzK/uoVB6s2tzOCImqZCITqCCtrWpjzZblNN7t/WErQxWCQLczex
botSZ/QzfHpt+p/VfhfyAuuZq6BvCqKka1hf+xiHHx+G/H/qp8wQhO5C/m2ysff0
FcWskfzE3TbsY0OxaP+AHC0ZoJ8klPiEEjajwSU6YjdfgTKSctxWoUoE1Z69840O
xl2Spx8DbBB0OHBEtervwX5+wMmFwbTEiiaNpe/tQsIRl8y8MReyeiyU+pmOVroA
Yql9yFWzZWhBSoz9dU/yf8p+N0ttuJ7I5m5nMiEWmn7WEd24JLU6f3+koWRhBedS
w0+61c2hpme4RZbklTH5koUvEMxfDs4t4v1zo486jUF6IWocRXUyS9l0azqgU7li
rLzqICYiCq/bhVhaduJX2AC5j7996yG+SRTOKlXRwWSIX5ueEj96oW3gaOkgg/Ck
MfU5oMbgsIUSir6G7r8yvToRKxh96X6d0IFxMDH6stg5hjR8wqQh2hmPxyGj2uUm
1Jw3Bdjpe8dKZvmCofv9YqjGYCwBw94dyXBT1HPUnqG5WOAUcT+xWadg0CZcVZxW
8N+ETcS4mY6W+3rFvuz8Dz2SXl/ou5Kr1HhCWlXvlRA3hwyBszyqWi/TSQI2UbOW
ijkTowWpJIM96UvxnnrVPpacQdahBBRAIes1u+tp1hS00OJnPL4UJihD1MAEeger
qJxVo33164iq5tM5p68XQj4JjefFx27sQkwTWO59hCd2tqqzkpcuby3tTsTub66p
pHe3RvB8XbAgahGcJlHJ57cSvvPEunqaNm3nn+2/V2sMNJz6TjmqymmnAOW5g2nL
76AV2ldtmjYu1jfzkJx2DL6B621+vVw3E+fLTS6pHRYUyDPmQwbSLC1uIgzn44qH
9QaePReCwnek6aLSz4d0d2Bew29XzP5iHvzTUsBXAmq7RurzOd6UK2LiDh9b9raq
oVWBDmjRMb35+hm36NBblwPa2KTe1wbZE5FQD8fkboaj4tBOtSp4RzLikb7nRYsj
DWKdmdb5Gib1swqdb15LPKKfbYWlyOnpp0QPF96JaUgOl0/xj5KODQ2zp2e6tENE
LLjJ29MuvNwberexXuUL3zOQMSsk1i29tQd59nHR1wpfiFki2M98JwmPY4J1K/OL
mbh2+Jfy+suyLuWtKDWkbL9oVbLhTbH2y4UGVJ8dxzJCCoBC5jGjDfbnrg4cUM2g
VE3Vz2slklgfRaKyad6zq/Bt+xcBIkA7hEPUi8bXPdXNaOdcFeTWGTLbFMZxaG51
5YfZR2uTSWArJpD37RdH6iwYiAwJlir6ls3j1tMgWc7QRwH5X1n6Gtt6mdA/74MR
nTThkhURb+iNIZaltWsKlSyXbjDa9nBo2DPOTVTOM72/o4krdmwPVHOlebyVB0w7
kTIHzsdB3dsTJs+Ft/dsnSWxWwNlZV8OC2sx0aEp/REtpo6hdkARNS2zwYl5Pgj0
S92oUTI1XL8WCO0teLhQH+zgKgzOFFCNCRcanxdaJeippP6a1UnELcJ48DEuQIse
RNlzrdoSyG9NCYPPPLxcU+INfqfdUEakzy41sgLWGlY+fZ3/bDawlmUnYbxlFs2E
vgTppN2ncHBzXGmIHZo05WNTxSHXJAX8IBaOn15E1QrIk/ZyI2jYvP48YdCenVll
rerV9b5J7O7bittV+4O9sWbxlvG9GGTryxvOEKPKXNiCxfO8vMkL8BhSDdVbjKo3
8+O6wawA2imOfGLK6NrhrZ30kf0Kn2L9gLS1WkY2Qje4vHwFL9o8bEJ2LzRXI668
ga9jFGC36Jy0LNFyht15wS5UY6GR7V6QSo7NPHMvXYmPIEMN/14zMBADDXrOQSSg
94VAQnOcn6tgn+XP7OP8PF1QF70JgHtT4Ku/HjjDtLPnlkKENltV725XuPfYxm+n
K+2tyzj/XQ6gNwIr9iOIpdflNvhZ7bOtTeYf1xa6RD2/hKC6yIqpvBk9FJ86mjJh
qiJhBiWiRm5Y0mnreTt8QKNpjZQhmX4hnjd4ULacTPyl5xQ+jFh7UjojRck2D8KH
tlf/tRtIT+d9Z1Yx7b3FVXJ041DKSEOHHf/NA0Mso8WCklXt7sSR6IYmJoby9qLu
oTdqEOjmlmsGUabUmEsLBkYGT8X2BGQP5p8MRI6jj4vEYtos4jVSK/yDX62Z2pr2
Umf6Qd0xb7HoavpkRLFs/oSmb6psqQ87OShWGP4xs5yNVsXMqDz8n5coSg6/6b9A
xX6VnOawbKv2MaEetNEoU3FAxwhVADZuTdUQ+GtJPb0CahQZKOKfuezDdhqOrZfW
Xr3q1ZVlEZrlp0aLG+zqspYlMkqsj5LFJsqiD3omJE5d3HPsgruj8pasqjXJz6tL
AceYXY+S3189HjhSu19nMf0WqkBqmCG5jG/ZJ1vkkn3o+jqyHfZW9VzmDjJvPVsY
865A/zCFX+pQ5EOJxvhps9miQ4ZzbhcfzBTWMPZxvSljRIpbMvNrSStqBdcG9d/s
269jSS4qB1FiqssfAovhKCA8hvEE0DL69W8hEqZn9u16Dmnj8s3H5ahmu6op+r/y
i4VVqZKprWscBT7ypLIvnhA0UoKRKyvjFGImUu15GGADAvu74djdHbAceUYQ8/gX
Yy1BlGHd1W6NmiDlIIIqZudLvQFhpnNOLsRx3WEOSbeXiqB+Wno+EHK1m2+ZNRKF
heLUTTK6BFVv8UVrmyNyYhU9wLd0oXeEELcPAg8TG9OwPt/KVyqNOxkirlet65/V
q8LH4YbD6qfNHxVujHlhAu3rlyKWhx9wIGpYZofEkfQjNfbmWVgviyMHBaBfRZp/
DhaYROEXp6mhwBIjYj8EmqCNfYwtMS6/P55dAiWuAa9yHFXCismTs8Wx6RzFEdda
cA5OfY93eakX7aoHXoH12k455F+mLSQocTJaeNmJiLMfLX90kuO6K3L8wGCdDlAP
2s7ESE8CT4ulQVZJWb8X4zwupg+LrlvZDA/g3OfrQzcOa1MalJRKZzBOJ+HIWpaL
t/p7lwNWM1j4KeW09veobyZC3wCDFQaMbBXvwjwG8hnXSW+sqH/ewCkSz5WCcqqY
Bz7UAA3bbMlVpuAvyeRotCS+3wuYSSgys2k1VETmVIXadrM5lMzyM9gNHdL1wkHM
4mdVKcj5zQKujO6zVQRmgFQfCTtov4EpEFKg6lG/4E0Rm5aaq20GmPIdOnmj0J4i
Qzvv5rzDBmA6Ake9/8WLacUmCIONM3gZGV0WAiDGhY2eOgH0gt6Vyj/sUuO8rll6
5s8tztylAHJW+ZNBx0IC7yHZHMw3gQFBlWQHxyQSgBBzmHl8cqvEcC2UCpNAm9UD
jcYM1pSK2uLDAKPt9w8xIKMDZ4fGhdavkJdQ2Z1qK/idbHaQtHLILc0HVP3FsWd7
w/G4cQR+pXWSPleAead/gTTAqb6UM4ZcGu4TBkX/8XPasF01STp6Z8wKlSMnkjs/
ans6BAKPMMISjuzVy9045CjCjNfgiO+jdIkQH1A33lpcUurxuXy000DCbPjuu3oo
oMPHAXUai28pfrfHHyAaBEG5xVutgeBrlFr72eebVxq8+nPd47yJneii/rO3GdIa
sObRLry701BLQR9A0WLbrWRJ/W8H6EZzMptJG+iPpMZ9cpcBnUNxwN9+PcX/2cpb
H1Yee9nVCdGaOw3zkg43Dd+s4mr8m9wi9tEJ0+5juH7BcfP4hyqVw9LrFOphc3eA
CBATBWuzWrDqnri5s0fgj/c+V3f9dxTQus+F1tUbD3aloM3I2K0fuuikgTkIzZWF
wNXQ2nz6KbD/iQ6alf3L9YvvorKLx7KtzjXCWicj6/XDqDUcDjusFOAixRXUBd4S
rC1HKeiHIGLRUUwy3IbKGcnE0+VT/DdEx7BiTZ7r2a4Cr4FQ8+jAiEE0IiEh9L9V
ywCEmlT8Ne4MLjABx0vO8dWXEAlvblggYLaYUDUD010xkZsiIEVth8uOT5LeJZ1x
jaIrZgnrfYAYnNGDruLbBz2s0TDMCV9x6YybyMWaxt1scO7UKQIUSgjr2p/wFvFI
Uljpyn+avCx1yP886d2RMXugtgr8IeTHX/Gwvwc8GDRQr03gXXTGVK2OCMlE85cE
ssrM8IO57u7AJUWGml8S9SHZT5zWGbQWeUoydLzbdEhJUSj2LaKQ7wM+MqmAb2EI
5BV368AE5YezWx5f+RrJ6ezHRfsi4OSTgFkbrb+lX3iOg1v2GOOAScMSyRycpKZq
7a1kRO56UmtJtvFSiQmZoCuLb/9smZitThNKX3tfwQ9hoNbOUpT6zhRCXFrZoAl+
sSZrl8dW1OlRDXIkV+kZkznw1vRN+gxlup++XKDBmx801c9eaRMt5tzWGf4m0Ohy
SyDzoHk6DQxTiMVHVLI5KtgOnnShmo41Xha14zAYWrTewBEPIMBSNM0lnb57A7UH
orwfjgvlLDi+D7sE/+IK9QKteqM/UFZR5dYvEXXZ913/AvTKOTd6i8eP1C+q5Bax
gx3Dv7xjKDhWYsj/ONAXFlAFEDJS3zYHTCd2AbfriI6b013G1WqvZ/a8LH/jRXa6
tWCBbpAmmGEyWoaiJuA8PKAqQaNfBGgk1O6e8+dDsNj5w5BjOOP9XMnT+N5I99B9
hnvfqhOofXV24kvIrOis+BeqoMJ6OWb09bmNLjQOmSRyqF4xknCF0WucrnwH/V9a
cEHfgRV0MVp4XOit+yhJfkSbgAQGavfW9gHL2rzE2G+XpPWv3tGfcUsSOGpouHA2
/B4n5SBx9mXItgFVouZScs7qPHQn6cefl5VejhoVlUIdU0+uYRuW8BPqE0wGGuao
VTAh9lxSrQgtES3h+2UML6DriS2oIuwhuX6muOblKTytEm8hY6n0Hddu4oFQ1I60
5ZC0SzQdvZrD4USua9Ff5J0w2348bCkeKgmagaMI7HyPq5iVZPTw5WbO8xoJfnTs
f8XXJCYkzTM2Kik51NDtbpTei4z8z5W2hxM2WJA75E4PskVhmuaQBxZl5ju0oRpf
vyL5ahaOpT/OuUxWc8ybf/AEe3+/I/axXayRj3aqj45/2/i7zIYwRc2q5zD1vKRf
HniNBB+ZqyIbiKcxnsoFLB/R1x2JJo1HRJC+9NJhyHUsR3ykQSAfQGlMbEMxHXkX
7pVNDVKvYsMrexMCbZUSL656AjEFtYDjza25n/vfU2Wr2EpW/Fhm5E89HmgbrrfV
3hwYAfwxMF/IaIypbeRtKk3Vz2+JBxCKD0AubUWmNPr5N9aaHYTPm0MU4JUvBQDa
sJhvw0rgdukoxzufxsul3jp/QKd+B3HNonnxKlz4y//tV6QL5F2L4yic74waloAc
BklHRy+gqSazte0KGRjO8FGwGDnJndgUYE+46sQdYtiVgl0Ov2GToNUQH2YPfRbV
sVOs0dxrzoUOizCgoyPOg+dVVmH9g1j/Ddq0MUuNnEt3EwI1CYPqnLzXjB28heLL
tRhoryPeX+clI2b/Daj1r1kJUuYrsQ9/AinD+En/wUqwrmiuyCuMA31osMIjwKG/
bInfzThh0wPnHkizvExXashFJbqFPixM6kKMLoB76vL3aQfy3YaA2N2s0kvVVuXl
KdexlYKw+Yw3v0PEvaUPWV0I6d72XeZY6Bki08QJNxei9c6Qxmtf+YaDiKlxlu/F
p+wQ2oAPvBKcRgC2IJSA7p2ngUmK821BGk/VcgbwIM4juESu4JHdkmtfIOzpEzFr
vcLwggvEIOYXEU8zuqoCOtaiHUTDMAsrAKTi0vL8Q0zvXqdHjCsYzTPcMK4riWmJ
j24FSpkpIeNN1TU9IgGEp4CCmtgKhYLVhgMiJylE/8jXWBJxxeiDkDjwrLPXW3u6
zTbuAy4GR/a6YIH2C4lXTwxB54gcjbVKK7ewmwuX8qoHDWTlzd7fcO6Ur/i0Pr7A
zyxAmdyKNIZkC9phWIvQZkmxrSdw28Quj/2iJtSWoYQgEeGc6bsILmYcOlOjyhtq
v9ipsa555XbktC/0iyP8wjhW8iwy9cXXUPI8TAbCRZ4iw+CY7FpXHAJO5HZEK1dB
Ja/u7qaF2HPokQMOEdM+FEVlA47N/lWzwCl83Engbe6zdaWYc5TqeTVprEgtIkHK
C/C/Pn8JuUuqm8UxkjbEmjnWtBNZdPAVknJAXMBBSE3rCEBXPTACbhXjrJd8sQ8z
tIRWZuPGGJMZ2L/g8IMGymsVXL1V5LzEdGfc8quA1fl0iau9no/D7fAuo4kjwwMi
+aAB/pXBXlB0uhpICFPf+hyrO+RVHbDhtTDIZCyZtt6lFk/H9xZuyim0DRbVTdci
vaSf1JU8k6rzix/eSN11GaxJmo/tFAF/HZgze1p+WgSeVGx0X0XtLDk3O7h2Cvh5
T4ZfJ7rwKNGq/VZbLv9kOc9iXBDYZW8usqShHLY2x7nIqghUWctUkLolDuWdBgEe
UxmG07x2g09SqUDgVci7rxpYvliy+tVYhtm+5iEPWBi8DYmVkEMhmCWoTLoEwYc2
FtJDUz9rOtwDIQnGOKlaN2/DH166qUUHhIBd295IKSi4n8fZlp1EoA7R9IbOS1jz
qsrhBfAxGvhVW/OePUhL0NYs10CJ/4tSHx4fLu4ML2RoeZTsXk1L5pGk8fGeFnor
JCcDGR/3uiyrbJunUwxCNT4ymSuy/aZ6IN/3cSL/am2WLdGxrcusP1p9NrC+MR2z
qV2g5lNCoEIhm9WqMFaOb/+qBpcUaMu3e8F9/nzZfQkGag1dKsK03knmW6ankxIu
lj4/0i3nbrME4Yh7MWd2WJJvh1sF38CpVukOer5J9WUJ4nGvH+T7OyNROIII28mr
icglzufey8sAA2hT+mxWo9CpxVN6kMrXJZPYuGw2p3qme84OYvX5PcTnNfeK4sUB
h+4Wg02sYVoF0ha+7ZJI+72ja0f2bkcblsQR95+ad+p8DCVav2u5zowtque6qm28
nUbWl49Sz/kmjJ5YJp4iDedecroAGir8j3PadsAHA58H0QZWnKoh1w5BMLbassFs
iP0tETV8DDBC4KrTBHdFYA5EWPsPSEm3DN2EegqkzT+HpkEL2WHtVevM/pnov0mt
o9YMwQC/GUONQy7ou4vVuFJ6jB5fNr780Eihvvy5Nwf6DTyfTLGRXTB+SfwtaNfl
juTQHgZObn+LSLux6hmMT+YRpnLwZuSz/zEhnA7V4fIBW5UEjcqmO0WY9/HjRzaO
xT7PaUh26RN/1800Zt577VOeCVA9gmXFf84+vUYWYEK8c2V6b77Y9amIYtX6la1/
yzjpi14+Mdam7eOP7CSW8KxCyxRj10TNwL5Mmi1uVCKzLNgD11GZySNUaKvQZXrS
OVSh+RE2vrh9FYEa6Q6+H/XbyLCRofpUtIFe2gyW5GRwjcJ9PuGkYePh/3Fsiqn3
I2/4wQhrsx3rdYj1oio2JINnpNxjyC3V6TcDq3GB/gRb3RrGXzld6mEVVhTwehC/
0EyvTDVyLK+VCk02Q9EKfNaHjqR2ZUSHtaRStlbX//tMNZosnC+J/pMiW8Imyxrc
nFNNnuzqEkFn75rfvqot65Y+hbGzi/J+eKfYrPcoznnebuSP/Ns8K4VaRREIZ94u
DJIH0R843vBjpo269+td7ST/zBqGn1RJ2ExlzHfKm3A2SCRnrfiv9SkycX1/OOYp
xSPxN8ooTfXMel2x9MrdgQhQhRns1i1Smc3gnWW9ABBbmub7YTjVv1WvUvg7JNAX
JxULQmSRqHqCnQ5GJ9YZ//5UfbACipK5BfGFD+e4kJ58Ky4eYSoe0Q9TIAMG+v3a
AecgD7RWfojlN30AmLDco+DsppIPpLixyrrD0c6h8qc1F0eGrX+R6p/7BdmrA1CF
SzAVdq+EzCUgtXtDYDg3qjmXoM0lCG4uCwacFwU1rbo4LAT8zfTuClNAc0621MBv
fXNPZ44uVksUWMHCUoeacahKgZBkODDFyDav5pAgw3+Uf6M/JTm39PMTaLwcJBKS
D0QzIKr1kPKEfpGluYzxhOVuExWSjTkF5kxYBoIhvnS/ogeNvdTKUUulb3c9tiOu
KCvd3Fqtp1305aK7jLlxigcv4Gm6EO0eB9tl08yMFlQiaPXEFOjP/X4HWEQb61XQ
rtr9hsjZRE+C2r91oy1X9umKNtUi0d1CiR9ObYi5iVKxlW9daIJeGwervx0qFHEx
ak9Cfcx/VpVoCkeWvy072qE95rHWgp1x6zJmLaAIBJjzXbRgMKlQW2eDiOKBjmne
KbsS2ESGj7qgczT87R+6qPvVHaLJeluEVsGGyM/LHptsDS56Oszm6IKm+OzpyBJL
kmUMyr1tURcdzasEAv0f0Q==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
e/tg5ovjyT4vXV1oBKFccBGokZQ/0cunTS6XEXp3YWQQ3jum3QJbDedqsd8rxlYX
6QTP3Nof/G4xGpLcZCJ8xZPCo7lf8Rfcz1QzdyT7B0ItAFcafiM8LEz3kezBdiV2
qUicx6O5EG0jUzKQCS4Owkbt5BVrsX05glszj4fSpsvarZ/NUkKv/nTh51JPj1S5
tgLlvTZrQS2PBn7VV9sloiWd5wSdztqfHqPjXLFa26kfB1Uc35v0H3TdH8DBPhva
gDrX+WrAO1rTkhcWHbEYJiTjXnQjX0MCtply+5zraOEHkHFQyv5qTL82JgDev7x0
/hypII38QfrXTBmjLZ21qA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5616 )
`pragma protect data_block
5D/FgughDcjhozmr243iHqh9chQnyrgfQzR+ZNu5Z7J6IZqIF/Y1U2ae5ER387i4
Mk4ojdJ0IrdEjxgH4PVPNMZSzao9eSNQ4nhIF48fZbJmzPmklEnjNdJgpRFtOzMx
YDnZ0bd09sEj40Odc0dKcSqNTanX5t/72Jp09V4dkUzjFKNrMmpI5gaTlI2n5CvH
qT7QF6LNAkiZuTnGGiAUWd8PCpwUb7RLMOC7oTXwDxMH0ds6y4Limh95YybDxuB5
ulzEhCXBmjVEyHp395D9rWOOWzq6TVCyHonA+qD6+EjvEfWbgKZOXG/UpOM/SL3N
hP/hktBcdlY8yVCc4sYJqUfRXocu1r9JGzEOQmz4xPdG5qfe+ez5ExMKSPvUOWer
tSxU0JFp80ALOdjKK6Iss3ZU/xaKIlLNLSTsd+9KUTN62BiWHO6S2r2XB7xQa60c
AoI7ytZQzhvBybNq2XQmlvr5PIfrJx9gnzpYbp0dIpSDfqu0eAQjrjsc1A9FrVVy
Vkuk05IqXZ72hLViZWuLSWahvjBZb+YZKPDOvx6uHYNQx2uJDXUEpAXb7xsbbNO0
RXMWN2ve45zdSrgPVojaeKZZD3dBS5zEUXJ9EVJAM403hrArkh9UgZpc3X02UJSu
TaVPmS4gIozmmB+tZUizippW6HHCrC7j0OZelG/R1ASDSK4fPFBZS6ae50VzblhF
8aGafnfTTqid/AibloPIb0j9TuaUiR4HynuJIlXgbjQgMnMjQy62YaPKDU1cDaxg
7atowqSI1HVUFE1uHfdkUkhb0J900PUOT/oLJ9muwFbMhHPYckn9Tkm9r8IcHxJm
EFAz6cT1ZIUa6eyUNEaszTpA1BzzkIkLUC43MLLlbQTQeH5OeGgO7byeKPO3oz/9
6iIXzTGsncINwaIJur/aZbyDXKGs1qyjIsW6e9dLG6NgQ0SBziHJXA75fhoXhoS4
iErFOFiB7rUAEZE1MabGUnTEUpSPd3Mth5spzIKQnS3isuZJF/Kpp1kX0kMv6J0q
2SveIR3cM2Md2rK+qfdA9S7vV3VjhDHXzk4y3BJXvspGFzpc+nRN5dZqWirx90PY
ewgqkpHChYnZaoukLF9/4+UouMGR/NF/5ov0RU41lF7hyYMQ4TpHD2Sw6mdlCleX
hW+Wd/HzpKDU6hC6rpZpvrD2rd2dWVMyCnQl5X/Ji4Rt6CPqtA9+p48RmjoYx+55
cWbBkhMv8n6vuMnYU14795bKMa6RSs6wETOIme+XlqAbuIDeDR+8vRlQBnLz4LVD
pbUbNFIv3JuslE8S08rQ5+WcUH3nd49EvawRFUjy+adrrHYZUzI/fur60RuPNzPF
x+pXhtqFgiwOIt3t7LDTC1YZ2PIQBsrlJTe0JCp6O7agzR5QFk+/OfvadBHMo+M5
nD6uhjA0DikoeBe2IC3qTFGX0nRn/DwcZDhIvTM7sBfFJESafLYzZym8WenG+iVD
EgGlsFRmP5h9rInQ6WXff6T1eOUdsrUHpavPDB7VFHJWUw1BvKDi8wjKk+qcRiYd
Kaw3FEJUmZn0b/oo56BFuGBPAED4Y40YY8t8mxBZ1zUvdcVkn8G233IevVn/SS3U
KiJso6tFTTlyVUfkhvDA7r2n5/nSZopTx9DWyCs+n8MsJQP5gryTWN2Pdqg+TCgU
WFTftgLLeJqgk7Fnl9xD2NmbFKe6mCb2zPFrkTigECnlvp4Frz3kZKRZiUyDAYs6
kmUJ9HR5bNWpwXNO94PmivkA79v78WYtyX1An2Pp75tzxT3PK/fBQn/g71jmMx6h
dxUZbt/Eh2Gy7UMwIJqt8LBg2UpjEB62TMokLcwKFNESXeKzv/yTJzJljxP4Fhxz
J3s6cqnlEFKbVT1wr6lLL3iQvV83tEzKDFcRBAo7KQSj9tWtbjmbznB7cLluan7j
118Pl9ZxWakAZagwq3q8ePecZcjkyeERsahS07SIvQKLPUQ+Y/l9WCRTmGXZKS4l
Ux7q60w+cuNn3UMC2QJvXPCNPpoPwF++9RhC3CcblSVUXRe3o4fjM2egDSB8zJBG
c5hNikARCusf6Vi8zLf5qORTd/L+IL/67MkOVag7i9vdOmQQmL3s2b05lW9wo5Di
OXAe15/x+tPhbkOkGHMe5EaAfCxbn73II5eQ2d6SxkMdYF7pVbsv+5OussteeUwR
g5wNVOaA0tGgjo9DoYydsYAfK83ifOn+8BIxxxkl05QcTkycXoxDYR3qBxvTrY6L
7tu/Ktq/4oJ/LuyA28UeYIFZPVOHnhlXGy1TZrr36I7iavLvaN77Rveh34hxkVCI
5rsoUm83/qpaceowY1HZgU0LEkXaG0TWQ7o8EePrw1qynZYNVhpNoek4JQPg2B4J
YNWAst+2L3qqnni3zHMVqJzxxXTYBfu9XQ6C1wrQ/lL6tcFIuCMRUUFy41y7ifis
4j3ihwAuCbziC6mJvoKcSVREQwMiaxgwDcd4oiZoydbs1ByQBrTgN+1u25LhAbVo
qculclzuuZA5e+KZ2SqHip6YZFElZuLDyqMsXCF3zTdMxrjNjM51FUZlrfN2AQyu
y85TVIwI+WZv7+sgdRgiUGppLNVBnanvilQA3ZIwii89QvKRim7BdGZ8+Shdi+oi
6nZJGPvlcAciooDjk3SHGuQNQqLazQkMFgwwUqxTy7sMdvf2C4TIjipFDeOf1YAG
3QLIpyqRQofmEseqvx1jn9sZjP/XXxtYtBHtZMAO9QQ8h3lXRFx+6w4wYYrWn9wK
wve10Gq02mq1XbKgmdiy+B2eJfFnnBDWZkIBUiCTKR8kjwTExU2cbEKmKjj/Xfee
wTjTpoR3gg2P2A543v8mD+bBGBKBFLZDv4YmUomrHvLX6o/qMtEvBof5zUddqpvI
ONxtpunEzKw9zenxQrM/odRl41PLSDmr6dJ85CF9K1t5LuZyt4qRN71EcHbsancI
uEWfy588ByF5DzLbLd69MEyrwsqQUdL9viQ6PG81+A/nXBzLft0oC5oxa1C0lNBD
SUoHy31+Mn7f63SeX9A2wu6komadzXzSjklkl6n68PoO5Vo/xq6OfulIfUlitllw
o27YPkSQ8cJcNTxby6XF9ECeZTIa9pZJxME31dspOoa6nm+uNw/ps3yEm93XDkMu
2gwH/ymWAAybXn1w9ldr3VXk2bXyBRTSNZnkEz2WuOmBffPN+DIt0gJ+D5zCayNe
5m1KHz9DN+oIxMscTo8qxCPmjYp2L1lQMAonWspmQrhe+2qD7soS9ffPH/2m5kxR
hoGTF9lkiCgAZhOG3xVhM6DKyj64mh5xjCDwjV/fpKR+lSXp7Deg5Rt/+3xYxgNg
KVI3vKSqzQTk4gYJAlnZVGbtKffKol34i/fdi+jhPWXxlNKCLJwdidNB9R/NPTKc
56jfXC23j4OLNS+HyZgvxenXoYY+G+DgW2eW+MU8eWg8U/gkxlxMPi+1gVt8hoS9
C9eBbXwPxX1SgvcmUIkOBf0F4p+8eop50GDV+X1Eu2QPQQfko41CNEwvhIXVhQpg
HTUmf198oK0vASKOdD6UgGQ7ZzFt2phxzSIfzyHJYg2NQFXuUkx35lTg2xA4lP1v
cE24FOmPvrGoWv5LTiIHpz78l01Bq9nnyVrQa/D3Y5AkYST0uTK2osWbw3iKAKC4
z+EkUMakaRyL2rUm7F393A7RXxUMyB+4OZ2Hz/jBCSIrqDlfu1OgwwOPnXOufCYT
oF9krK5m63kkPr6YpRI2euyJuoV/yqDuioye4QtwBIe0FACi1BE9Yxv5Hg/J4bh4
YEs4S3l01NEDjGB9cQum4gQkw47ohjTG01wVqpARH1fLAsr5SXTp/VBCAV7/8sCd
yX0NOCXz8NFlGtGBYe0eX5Dub+2UNsBY78o72UZFywYMpamSKyONHFOU4TWa4qq7
1fYXJYX316jP99BxFc4hAKP7vq/4g0sBITq+Ge8TYgVJQ3tIqB98dzoFEDE8GXG/
J/XKMHs2dJO5SHYcQcjEUed2MnoxE6Bp1W0ueDUUNAd/jECARvKuAcfbspKSCFlg
vCnJBkM5MBJAGGmRdlQCgcjodlkH0sGGDbWVL3vAeOXB+8nM6inXU7RdyPozzyoQ
IB6rcq9QDR1WdtRFLmB7WO6+C4mw55IcEhN2i6mzs8r9/aSA+ZQDwnYHsxM5Ow0l
WgmCkINX0k0dJGMDl47DgmuMJ50t0sbCZE3oMN2x0EMHZedAfjzy3CK6J2GE4XHw
WnjDINuKbo2NycI3X5pw0tGsnkQjRY7OZkmoxRGOys5UJ87z+g3FtmC3AV7L/JMb
iKp4RtlrvebL4low87n/ow6BfQh1Fui4XNQiIoAeNd83aTh+HEuPqDEADfuoZQ6d
7Y2UOY+wXbMrKwSin9CkZDWXEhPdW+eCA354ZqLK8jXFg3y6iLHUwd3gihPR0MeM
3Z1d+1lNCtunCyhKZVG70VhfhE9MHUz+4jumju0XDAPWt2cxV6LwXeu8aBPMqBc1
99pb1/NY0Ldo6TXZi0DAHdRc8nLT2wo4hFYe0Sm54h1yeRqYHJ28Ft3RXWSmMYHQ
h8oDZ/23JU4q3TfSiCw11HmcFfKuHmPrltdcBLgh5LOG73ai34FZCYzJ8BRbAuib
Y8hAYkYzo9CPrvVBIQPrLJtlL0u1SPeRSLyU1K8WWQUqQ0a+8hyHZW02o9tyJIdJ
gmtWE7gxyeiYbhg73Bdy4I+XIdpDXxJLCCcX/os89aMbDwOhq/OZJCW8pk0EqWgh
XqSaodUSY1vQUW26iPdagKsVP4W60g8Kc9zOx7M8vZP8hXJiJMzL+jEGC3CAqBgi
IeHlm+Kc4XJ06hIZjRouVgqeDdEoS5hTXZpkaw3SoxZ+DGPZfCpKiLEVkHYevh8Y
OX5LAcaCEqtZm56pbB30ZiANyBmw344LI4YsXTyFQa4Xzif80Ak6yfu0youc9eA8
i7rGFD/YuBh0E+5D3xBopGKm1/Yclx/+Sx1HTRqGm8ZDoZSkU6jmZV/XS7IJItyK
baEhmrMd31lwczA0ZMaTshIfv8PsYSrM+htZ6aCXexzFvYaj+q4UsqlHVXVQaaYx
UXi8D/bfL1nH+kpfUYeTr1NVlZzvHgaY7AbkerSrSw5wmDdViizV7tCYpCvQjhx6
LGC7UcPHpi7UaGDE2/RbThqpzbUBjNcZLWKO19H3mslGtzoajZRM/OKaYz12GYyO
ISuyTyQq3tPeVwvg7Rnu62pQyJQmgI01abh0OaA0imvS9Yv3AiBgcK4dd+GLOk8i
rjmvmsSx6mVbYC+L3MoeqG3kh6G0yuaM/YkyCLbegrMNcCQQwf1EUC5iEqknghjE
SRO0clbr/yO+zqaM+YPTG5WPtWnBGj5G93boeAUaWZOpCECtKF91cQGDs+NFOLAM
AQ6+4qGgxAWkPccONY8fymYcGmmn8dAkJnwc4bJdIw7VYiycU2oUY1EfdGRczzz9
b1mln9jz1QVlm+lS2WG5EbUQMWabjcvUuZkA8an9P9Z0fzGy7gPD+kGzc/ztNCOK
PqHpGLnTVQN1QWt6Gufsk96Zl0tWkOnHzly4W9Z4Vd35+S+OS3nE1VOCg4Bzlfge
tMBr+Sf6iY0OV55oFFifsz0DU6MeCgF5fLPXVQzS6wXz6fnZKLlw3C98s91VFUQD
4QwWD11ZqUWyWmvgZrSThsGnUZf7fqu8vbB7OqQ8W5yIOKjAFWsEEncnZ3Wz2tBt
ZpURx+glvtgPCtKNQGANtuiIcvMMU3LcQQT539xz72hbQSmZ5+WBZdb7S+OM1nOw
vRJMTVs2qEV9GL3MYXnl9Q3Eyx8nNjRKayfKDHF8WHyd3FBs1ng1wKi80mE54Ilw
7yyGAmxw/VuFSftrywC/9bPyuqIU2GPOsxgZEqIin+wSyVlsa5PEeO0wBrFk3TxC
q7lZmR57QOOtLkbJZuQDo5eDhYeqH/6llpI66CJzWH6SxuIcExUYTHjZKerGEjxa
A5OT/KQTplZeInzehqxX/YBEW5gTYi8VIBq2DYp0VKTFK0Rw+3E8xUMPTkto7In+
Dq/48nSy+rApbmz9da6vYixhJ3tPljs5w6vMuwskhLvseUpIyBUOW15bVZAcMwkR
x4nHZGA4kXFWMvusit58LuVf3xqIi3xRiJ4CZEba3tAXmhbY2vlqk2llqG8PAPp9
2KyeuZHzA2khraW/hSi6q6VVlRdpej/OzTnOLxtTaF42vF+0lIaSOiN4iaf2HBmk
HPuUuQtpDifwg+S9eUg7ywDVvIBwY361h+qcW1++mLhgjRtpNALHjd93oZA3MIIW
xLLQEnBSM1CVzH/QFYUl6KuLouYmz+Gpp29lN3Xqf3jKgmxvcd7osK5rXHdTSlaM
wZB8g1iNOXFQrvgVFx0qIwbKFVjUS6Tf7EPeDGGYKn09kLVG/BdoRw1eni71jRMu
H2aTk0g6r+U3wesmDh+0EsycE7+a8ExZg5vJ1wRLDbktasdA5E53Lve6IH/N1SJB
0v8stlz7gSn8Dm1vuSH/fwhOVhsS6R8mz+vwP/Ye41a9y06pUBEWnE+DFuWUHsFv
uU773ejkSjZr4h1NwC/THXsJYerUR8fWsxbk/rdO4IobZ3nkpNLxgCgy7G3RzRl5
xplN6GVeIzY/bPmTFrwLVRia+eAA1VHH8Vr6Cj5ix1C400ZnFJkwppqattto9mg7
iFhTGqGGyXjj3AjX0BUoV6ieLLtyZkOSPhQraqOjgqf12seL9CTBEC6SVz+Ijlgp
A8IGfYq7IawA//qILMb5igZKZd37ObSGJ4SR+qevM5q+PToc+km29m6iA2upzYD9
DC9oTLR0D9+kjLTw0jgFwfNScsd0sF3mSlqD+t/+0HPm0VelhdXKyEewKXRMR9m5
L5aE0Jb+RGX/cIaVzpv+yp1rY8y9CtNawYRKUdsPwFzovW1DZove667FQ/Q6s2h7
DbEk4U8PPN5wpcp4T0Yd8elJ8XTDdnkwkgTf+CFppa2o6YedAjJZ9fIwalcTrKkB
egcyT5z9rbLSy0YnkLP2PbrdLz4PfSIgzDip0QQoFhk3uYnVj5uCg9ITv3JB312O
oje23Yfr/pjekUHVg4xUpNzs22UxuOGXyU/F5v/UBfYPkZl4nXfx3G2lAEG9KMvM
C09I/YKYlVcBjpYSKCxA2eYg1umGmGQKnf6KMajXST044mpFoi6FZB3MAME56v54
J/2ZTqXu7LVX7k6IOmvkjzXMUQoRTv/DUbtcmEhbZ6UJBhgI1D71upSUTBFx7SJc
LPcJKfMUVzG6FRvuQDAiD11zgPvgWF/aNoQgFdW15WW9Y6IlXVxkc08I2Hp/4FuP
oPOTn0VIdQ+jCugYT/hiErXC73SqvsnKvEtxnCn0oMaT/TI1fVGXFa17HI4zjXZz
Q53bc7Quge5n84BJKQGoAjFZVdtA4VeGOzY1KxXTP5Z7MC5SvldNCzesZzqt9XJj
393WlRzrWAZWwUotMYEodpZQZE3MEVxrZJsYmhlNToxQh0GQyZWBqJM69s+Aajo6
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
g0SvcjVV7hkLSbwEFnNBoPLpdf3dT5q3JHIFfSnCoJaVGKT4LoImZ2Ewe975Erd3
IDNNsNiKAOy6bocLQZ9+iT5uR4MMFOu2Y2aIbTtWShRGPiLVcOPCxPKNPi6E2Hcb
W1NNQtk7hu8YAthUJzBT6xO5ng60GJAPrQGo/KUVO7GHwLc9JtvCO1NXPCgPzUFn
TfZpZJTeYzQVvW0WtZpQdrBOk/BXKrJbGQtbXDAD8XgGrd0M+3T1czNseOf5WISi
ubtwHYgIo8IDJo+TRH2EcB6lmoMqJpJpapF41hGccSIa6ICksYNwJ+99fh17WXEi
SXMbnnKePRUJGHg8em1d/w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6160 )
`pragma protect data_block
+vX9mvzOCX/Oe75+gkLi1Sgd/qlsTQyi1s6Qc9IngZQJ5KCDO8a6dmbZmK2JW60O
LylOzHJSGtcAKfNdyuLeP4ez9qK/erc7ehkBacCJXjk4B0FrbJzRMJuVquIr9Edx
Ene60iAceys+cMjtJ6wZ4KoMFdnM15Uhl1y0ATyEsX1k3D5/vwVJrU36wuoyw76T
uPfaLm3B/A8BKm3kStsKCmA+xa1q6CM9w8Z7a53VLwSOCdzPN4txEpOIbs8URJhd
qHvHYof1EF1gfr6m/5WYvL+AIBIpiEA02yVqAHoPLS1U//AdUpUaoA3YcW0P5Fxo
1QZ797siSrOx3HrSxYMhuvH+9Njq54eTtsxy5jBu1V/JkRJ9Ke3qa1Q/aB31gmQF
syGkfI+sOi5UU4jpD4CCf4goYw0Ed/onC0CJQu+74QnOIuRDPGDMVvZaEU7Lu913
voY7hdgXV3MunZTAsDToScYGgg9IgWQtCOCerdL7GVB3MfTq+JJ7qMSWy/jNbaNF
W98dWg2xRyYeGCdcBc2ig3bKzq8gEFeaKcf6rtlHwugCcHsiRwxI3QT4udxtsmJL
UHuppPUZpc2hXG/G0D5Yp3v4gbEc1EXQVT6iNPg9s2J2H4p1eJSwwgVCcsgbp1Yn
xRMUnm/I9SXfO+Z/VlVYbzs04Ww/JXJtguQpurFqyI7F3fabEJf5/+UOEnreHXUO
ThrPB2OX/kGLvhUVjGFSYo0lno7NvRI+2X+DJ4voqTXDXkrnCmhS9t0PnHH9wgcP
j+qvhmxIRsFekseRQWgS6lbgNP2kbVhVE+GLcryTa81CZxunEGj/eSV9al8XNgRZ
7+aDbk5NR9ZRjQmba+8F8Mir6wwqoOJpcwjdKFgX3CQxH1eB01YGkgs3QRqnU1PZ
qvVNiAb+jS6yUhpD1znh1kjPQYBUk/9EU7s4EEJHhB8HNZOc1hKbITgw6Jx8h5mk
zbVf0WJ9+0KtsPEDid6SSMxDxFj+NKDnWKu1bAvRUNko7fGQ3h1u0qubHVZUuPzu
bMOM5FrOMxrhUaDGXOQuUe+nNX+iVhHIBmOhq/15D2HbIcXvNLiXPrHf/Q1ihEUR
g7VBGKMuFzYGhWJev1jVwTyTjLUg1gJy3cT34cgiOKZJg8FKy0aLP3C/p7RCQtz+
WPvB8mPbeGNa9x8h9X0+ce3uB3R0dzneXOcr4EFziZoRh27oWZmSbubYrPGpn2Og
Y/TrZS9L0MG9Pu/YHjFki65zTplZVMoG8SkUoxlYvKxpMttYQml2hdCLge2X3DH2
q8p8uLeMDHlhA6ONqfXdyKSc8Jgf9k7QOKjXdqoelxAbLrmTaB0Ww3+hbzOibkCU
sQNEew8SZpHSo3pim9lQdP/uXxgtHslrnYweK8kgHM40JnIKxjH/2tEV5i5MpMCd
EAiX6RuStbYyUA/3k/LUwtT0EV2Ud3AxcVZsApRTBalKd83JTVmDhp+/yxmA+wAA
nu6d7qyv2UdNWedcrwwl8pcbrmnLMQy/W69b912A+IWxQ4r4mXz+eZ4Q8nAU5gRF
W4EQzThdawrzQz2mLmr+j8tcdTEWWjgcKXhP1b+nyCknK53phKUaPZDmZKcJN0Ar
PopUFwJm1lzU4xVpVNxpIMz9msoAsBdrLzS8WOmdJMdtkUH7INNVSELLj58evuEH
CKb9l2Zwow82YyFhA91Q9PFgpVEK4pm6ovcjJma8OPPSbENbr0iSIQP3WIR5nKvt
mFUos4nOuiqubc3DHHA44um/aq/n04e/lc/HUzJFBR6QNkmav+C7lRy/d3jI8qbL
QElwY/xHFzA4cZYm9mq1qPOdlPHcXZyYFSTTu0KgE1WCMjvPIf4HY1BxU6aZEdqb
1aq8kFZenLuak6cwF8F+bwNnFV90X2hA0OJFEfOSRhJrnu+56Aq8zeJHtp05qpe2
2tWqCqNjYkYonL2pDmlfkPJ1kvjkqzgODgVgQWdwH2UwBnCCEIEZ9k0OIjA52GYc
hQNmyUiXR8SBbWGEI65sTNOTttEqb79TLH9vDkrJZpK+3UoAnODgVGSdVM1yqxZY
kCXmwsiTVPX3AiGhOKRxOZjmneezR5HHLd78EFBvL6drGG53xuI4VLaQcSQHI+Gp
6ZF5b6IfjvjuWoDlqQ8Oqb+THWGFFZqQq9QjDTG0wZ58aX2JLVE2rsFHZqDlY04C
GT38XkN67hIXuIR3Htp/r6peFi5sz2EDsrEVd5qNowDRhMqqmg48TAuqxGrqTeGW
ePa9nygO5NyZJeS3KHqBTrC+IODqROG9aW87C/wVa1wE/1MVr9eWq76xAa+PXEaV
s/pYgkj9fN0NfL6XbPel5JzZssfJlRtEsKn4AGkm91vaWv0RBChGNwxXyuvWaXLj
xV3gVkWgpMsChmp/1V1T3PeBLHl0k6DCaWAbfSOGaAETmGjkGHgNq+X0Za52Bpzh
FSYIc4ihhdZqE5xICNXN/2xfCpqgUA61mPbEqbulSqt4O8sk6Mbb4BykRp1z6ue4
23Y0Ws5zPRyClBMFAFb4R5f8TBHJLbePtT79VvKeaaXuZKRAhCl5fE+n2CP4rHNY
ucVL3MwmPUtkmmIjhA1A/xY6ozUO0K/xjhaxG8CkWU1iwhMuO3Qq/5TGvKjwRMz1
5aBUXlywbitTfnzGiJUVAKTYThxmEtFqXlzxuwHDJgjl+mJonbEtt9+xRgS4Pi3d
JcK5APPEPBYA6KGmWEU84X1ovx+Yg6Da6bw4vGBFeYsHQUd7qMx0VTYrPtwoOHVj
O/C88K8OEaUYJ2e2kXlK6O9RL5tHUVpBPpYtqUHslSB1ApwYRc6TV0uaMFpuhAI/
PaAa5nflUDibSAKoDNLYfzg8XdslDHZpUxckX693a0ei5DRTQSbZsMoQnXBnYf14
9dpnpBYUSq36iQHCtGiUnKFfN5izkDPxpMSvVjpK4c6ocFTCIsG7ZtInwOYmh2Te
6/r8n0ERu3VO8Dwm0puVrmicCh/MwxV2FALwYxRWaoT23kncvmxrIxRvzVCjDm7Z
EruW+yMAWAkcLrhtOnb/UUgVl468+bgE6xbtgFsL/H5Wssb+wCvcH+b2ARhTUBjM
EuKIg9XSTckgMLLNWULWxjXCWVFteT3vxsROV/0Zi8YO+4iLkjdpJKEtdyVVG5Wm
4zXdp/ozP5IUFXKQDr1Ox8+Gad3OZNWOcFxWmctMBlODKtfxDN1MQQ0un5ztGJj2
uXRqehbHZRb/u4u73/zPXamS7QnSqpMV8mUQJh7URDO9Jt/o4wIePcgAdLh2C5z4
e+6AefRmEC182K8A2Ve0WSdqtnvUX/jci31Tiz+T1tF+4F0JYx1WatWadWJH7FHe
Tjbc0fFcdRTRHes8cQ1vr41h2t5nxmVeevCdYpw5YHbXIGIySRyxyvC97D4K6Awl
ytCIP2IPxOmiTLAyDfxXmZeoCWM1XR5occOD0O5AqkbCHr+NnHN5Z3TIu6+wBWzZ
WMCybdWFUpNg2P+YQVJZEcCHawFpFMuZxu0vQEJws6yM43Muy1pXiDvC2BoVy//k
ytkS++pp9eqgVBpSbj3IFdlattViqIlcRYOmrslqglYhnNeauVvaGDXKDgBXHKlj
YpyTeA5LnX8gmgGcrSTgmZn+QFctKNGxWP33jmM+mP2qpG0AjD5Fb8Ob70fVXaiB
AfNY/ZSI3fhupDY75UvkNchcn4r+trMR3WP0wt1gcuBRHLqI9zLYCpayhdjMghxG
FWArh4ik6Cw9qrDtpveNYPTHTjL3x1cWRypwGew/jzQ+u7U41YeOfQPtyIFOMOTK
bfrJOzb7UjVupYfRmAKaopL+9Cp5D39T8ryp3g4HcTnuhFBF4nxIE15SwIuFiowI
L/+FSg+sBeuuP36dWyQh9EamlwCDCTRxhAOQ/4y9EW5kpYF7WEqc6atqILXI1Fg6
6qs8z09Nv4pittymUk0Lc7+CqHe5lgY9E1wZrguCgO/RzFB1DDsXcyMx8G+/Kp8J
4lJthzDHwaiAln+EM7xWIwlBYhun5+ZuusipPpzN6n6vX5jG0QMDtRybvfs6AhA6
EcUmtC5vPV18qJaT2B3suVxFiQBG1wNFH5HIVuqbm1AW/mchrxBqOhXF2nWv7tN4
GdVPngLl5vvuFDC77ozfe44neDDUdrqrP6sdaRKoZ3YEfUMIbFtu1MVCEh2oB7m3
YchFl6CuDANIdz0BppXy5Kz3G2zJDzmsy+WVYILYM5UHfLafrNtDm5B7XKR8Ax7O
/aTyp/N271rPCMNuje3dQyXrLmw/zYs6Klc4tp8ZS0/Is3ZSUvxwPM+gq4UA9Irr
n+SENZLGkIgW6pzdlwNR9F3wt+GEuuy6SM3LvevLAuzz235BPNwB/0lJ3U2Ldrna
chf+RMg+LixekAS/dW+2roopy7iE1uuasOEJidFy9lQn/6gj8UN9x/WbqSyz7MYX
XvviaT/mPv2w0BhJQD/hQ7IPrWUu8YwlH7LTsOCVYDbyDV/3a+O78C6DzD/wsdYR
J19UUw9nUZ23uFo20j8G/9V4zTVh7Sb9VkQXrEMORU5OgElyn7gD4F/IEobTlqhv
VctoI7Pw56XVypdwrQeCFYZp5ssmWtoVTN2X5MXV5A0Mne4TGzgmEnQ7xH+5yKOe
IYT9b96vbA72CrO/tWdNh0tfhoAhogoER/olnIEEhk8RXqqwS9NAJd+6ywHJnMcb
TFp6cY4UODds1GWbS5M2nShWdsLS1NqyEsHgTp50+pBaSqgQrAl5cp0ec4p0uDpY
D8iOovpEBWhXNoLcfzcpVBMDVlrE2bVLu0sCO5gCmKgdW+ENw3OPV4EYn1iCxpiA
EGeC/TF1Arm6qMttDhR0gSDxdTsXR9mdiwF+HJk/Ki0x3l5ArSKfWVWwgptcn4Mi
O8jwB7OayVsWB1fPTAAhDHZmOO1ch/hDYAWxPlj1KQ7JS0Wkk0gDZXGzAiHKF6Jo
9md7tTZHKN6KumN8gPCKrFq9INCvAovic0pChGZj+A6gv2I5yn49RYUuXbBPz7Xr
4P2PRAli4cHp8qIcw/yYMbXIJ8KviJEfWEAAhRLoqh9f6hVcyuKS/gFu3axOf6FQ
llLQ2r3WNK5bfly1w162N+kVZYpTI+7ZG9v91rTJHQ6Nha9fewXDwVla0OxZcbls
LLrNqx9sxtIoj6f+zCtorgyaMEPn7YKP/gMEacfbEcyw7b+3hvFFVAOWVDrm22Ib
vpzaHorfEptkg92bVYX2CCJtKUSlxIYwusNOzjsVt2vN/rrV4lOQ9WMtDY2EsdRl
ZZmhRhdJMyRkuysjv5AF2yrGKiGxzkR1Ym5LXjht02BaxQ7JmhWqawkvDBBvGBg8
24EObghH2ple2vDVVvNWkE199YSYhiHYef4cv6m6kexmb+K12dDLrH6LOCuJOgrR
YtlWw1EHNBGVVO2+BgzL7dNXpkowz+EotN/0Sc7bsIEoySTG11p0U9C4BqcxOOKg
JSWF3dHaFndYUSu0wjgmJoECU1Ex8uRQp1YgRKRbkddvyyTmdg5MR2GVoeoXxcZD
k7yas8BSvnAnpjEqeE48T0oud0Lvyhh/+o894K6f/8V4z+rjsXVuODzPB81iU9GY
JRxrH8vumnbsAHR0qsasBJZq8k2irTzKv+20vHpf7tsN3LKmBzpLyk/cjpLplOv4
6C+4hk5Kzt7ehC3wQh6vFOTadvXh+AMx7hiDENT7R5gosoQ4MctZo2RfxN/7Lc02
ZrETENQHG75Xi6oftdaL+RzThVeaiDLJHbhHCIoHz96vTDgNkEiqOTacX8f27fBr
sWS2Q7Ji2uL+gdoheNYpALhRT3oqBie33SUeBUEilYLf+0WNP65oKkPoivbVYNNN
i/ACrFVbAS/DDLDlHIRCnrlQUcVscUV+BH9TbokGE/FNjJdhl0yRHlVAhoc9Y0y/
78LZdu5h52QP1r65PAGdcleAxkwfKKcWph6GSDkDT4TR1a/4Dg5x15mrjLNbdTtX
PdQ2I7cDHqbLppjsCExcHHObTUrdjy4DjV3WjcyiYVVFrOCbwHQziToUbimDaDPS
DWEFPS2d7weIFgI172Wntk587Xs6sdKMQstJU47CwsDY6NC/R9wqTjIk+xwL/saJ
Sr5YvNLnxCJxWmjsvHT+w5qkJiyUim8xGovJkhutreAu1cNg0tkrydmGOd+NwDVm
kCXxKi55AtNfKbfnOaQNr2Ru0lUqyrJZT4D/K20djBrxnqnSfjCwtX4BgwDVWpCx
ia8RG7DOnq3e9pB2HMLpSYRdZDaqvjt2MCoQQuu7v60LQqVmgb9qdj4Eb0JMpZwz
+j6QRDpaFUmm2euknKN6zvKMmpCEkpXBH1eLaaARSOhl/mhsmrasOtbwET4v4bFB
C0SoMqBhG0BQlTWN5GMgkW9agdIQe8KuM9ul3mJPvMxxZ0REB4pA1gjpLBEtM59f
cawSZ0chkQda7G64lvQVns1NjS7LkY8jqF+3SAiIRqIvPCWSOzeFJjHeqiGwddxP
uepSWcyKYLKd0Y2K+Vor/d+JPgdy3MsaSKRabUzGjHRdPanAHFXjgxrjRfuzWmSN
/T7wNErVFmjPz6+4Ed1Co4q4LCQp5kbA/ZfhcKpxV5Ja0Wuf31jBcebpeVq/4WHS
/jhtniZxwefYxWnfxzBFfqL/G7ewcK4KTubidhJSd2bKLw1Ye4CgSXAvVxmOtM+M
8o4vYHDZHJvmo7VTBkV3gr4oc4maXT46fNUIoSYUKIYRQ/XUe/ZooFpQ/qMuW8OX
56RwOvWcnuKcbQLOfoc5Q6cZ9MGkV4Vzmk+Df+qBrjMx3DNxdriKgygxkB6CKaxX
2wmxFR9XnouPZVHHaUHunLH2j1HzFedepXmcCQHcn3Bu6r5h37Htmcm6yMTB4Xpk
Oh37Q6r6FFIB37H4KZQnZRoH/V8IrsMzuZLV11GtrT/1K/tUEQrrj4WVw3QsgHCj
mvwOgIH9C9KkgEv+ysL12Wpxb5LLkNwLYeY9TgL+4+CKn21wp35HqxJj76dxL0Zh
MYneuIBARNliURGC/t0FNjo2w972yluL0CShIEmRpal9tPXAA7nYpzd/49dtZQ4n
j0VrJrBuAa3stRfvVL/vTnDkGl06VQuwHbNQgqWPS3oimikxy2nZGwRnWDEyhRx/
Z+2NFukWhY23zCSxfm9aEFClXoNe6uN9Yx5MGJ6QFYfBTa3MDJ2oriv8rD4uPabR
phFO/pyLok2KXdOq6y1iVYGhbas7ZQu5ru5jOPsggu/oojBvm3Kg6J1wqRMhLyNJ
3BRVQihWuJRhfIIPgZDUHd71qHe7QAElzqo+iIEM4zcNqnO7OVXDgsXDkGk5cXVf
sEd9vOIdO9ryMtB0F0SUcuBS4RS3xn6tkQ5Dh+52O8Rzh9Qd5UefcLib8mf9N/HK
AcyGHU2mvXV6EceohXW1HoDQL+844INcafKW0snotfuP5EYRudYz0khXJ2n9rS/w
ZM5RFBSdUIzoSNDH7331JhJXLrGaMw9McgcTRJr6+QHtf4NYf19Pc7e9FrUnR+bk
v4HUd73qEtNtEPtDH06fcE/6ux8XlMM9dQsnXRHz9Sq3umz1S9mXiTTUin+ZK9W3
z11jpKl7n2xspwzCLeCCtvBr4frDwUPVlHLuW1eDjP0PodNMY9Isf0xDvbaB5E+1
DB75nEUKnwXMmMqINbeoT4T+mLSWMPNCifWckqN/pypEIU55imST4DGr7zgZMCbW
/oBRhxswaIkcKiSJFjDFq56HhaCG+VQOD9W5iXZrjo8AsEVFGpNaRzjsf+FMr1/E
vh4z0lZ5DLmQGf/RmaZCyTOnF2/iVxRsI5QUttA9sEDY/6UCQOGwalESWhzUsSmg
QSi/SjpLICNlTRGv9WLJU1P+qc5iTr3LAH7wMOyARUOPJ6wtwBtKMICXJC4XhxvT
0HZDXhkvyMbJdOz2vj73lLCq4jWmRI63POk+Z0pB5o6NZUDP5J/LRVt4/d79m3mE
SIiE2gPBorphssIPGTaSYJHrZrDbqWgyPgnjbRSP9w59x1/hC+dsoVQI7Ad5TTXi
9sMLM5uLAzX8tghM9pqtxaoSrG1DXTZnGyJOKtiZhoCxJ5bZw/HklIhUHObHw1Sg
Hc8+RWia0S4QgK3gEG7y+slkrC40xNFAQuwNgXQRETLQzKLpp2211KtmFtY5Sv5X
OppGlppgcBVgt3oVBBJWTzG9NTgshT7DIF0j4IL+ED0Y+VHfP/xDfC30BwNqg/ew
z7cj2zbmwz4WcjLoMgBrpg==
`pragma protect end_protected

//pragma protect end

// synopsys translate_off
`timescale 1 ns / 1 ps													
// synopsys translate_on

module `IP_MODULE_NAME(efx_asyncreg) #(
    parameter ASYNC_STAGE = 2,
    parameter WIDTH = 4,
    parameter ACTIVE_LOW = 1, // 0 - Active high reset, 1 - Active low reset
    parameter RST_VALUE = 0,
    parameter OFF_ASSERTION = 0 // 1 = Turn off PULSE_WIDTH_CHK assertion for a particular instance 
) (
    input  wire             clk,
    input  wire             reset_n,
    input  wire [WIDTH-1:0] d_i,
    output wire [WIDTH-1:0] d_o
);











`pragma protect begin_protected
`pragma protect version = 1
`pragma protect author = "author-a" , author_info = "author-a-details"
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.4"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
n9GXfY6k/ZhtJD9kiUNVLtaH0OSdANAy0snKnBtVVWQ6QOE+Ndo/VTZDI+hGg8g9
BQuVUO9VYpfcYCQvBCADNQKgSAqxFZjzIRV27HIOeZCFcQqQWxv7S+5zWngR1OAV
+Gybs11Q3LoZ/IBIGBpd0XnkdyubJyu4oBd3pKxGDxxRxImpbWTGclPoIrWLQbHy
BHYzpKNiI06B7YEvoi3X/d1pKZDVylZEMUSddSlug+uFiiaJtWQh6NA+z/owDEDE
V6bVUxyNm5aGjXjEzEECUcMJcfeV956Wj1jl3fVxGiNP0REOhvPr0bI/Girb6uQV
p+McpZkCfrqzEUBv+tF25w==
`pragma protect key_keyowner = "Cadence Design Systems." , key_keyname = "CDS_RSA_KEY_VER_2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ANz2D8YrxkPjLNtSoqQ0qL/n/jE0iquIWk/3e3vE+oIaj29rVvK4slX1wAMRUX9N
upY9Ha7G82YH6HOWpzJQwnJ2DAY0Z3VQ3OFLkDk/Huz3SCQACFeCg8JTJ+gkqyIY
3qkzAdDWdipMtrWdFBeESV7jsaxlunckrpbgbEzci0JaAN21i098RIWuzrZr1HTH
dhLLzlbWTgr2KnB5l9x0HVdJAN9fzTDmnCmAJMU6tkoHiQaAhQNuBUDo0LAEd86e
FLJDJhF15fh4yrlIrzYr3WEqxNEjnYmgMEPuSLo8lQrcsVIomt1zamkCO09pKhfp
/GUCfdkRxv3JWfTNRFn7gg==
`pragma protect key_keyowner = "Synopsys" , key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`pragma protect key_block
Zr7q0eHhaH7ptNB2EeBR/IQwCwGbZ8h5GSZSb4880yuCpqV3mF4LyVsWhgP/s+oL
K0Ls94YLsw+5IXRtW0LZarLJwXt3vd7exEKa2b4yrwhA3xkg4lvSFlzHYvUrejVb
pvELZpNMkl7gKvWAY1rITa8iFy4DIl/v0EZIF0sNnts=
`pragma protect key_keyowner = "Aldec" , key_keyname = "ALDEC15_001"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FuzzgfHyzdkm19HzCmIN77AO/gXQ89jPquRQ3E29Wuyahb8Rb3IaHBb2xF+ucNQz
iriPZJpxHjpFDU1ldMRZs9rmKQ1IEUkfM7Uriu9aXykiHujm16In9i6+P1J+GMdX
fZceSO0vZqr7OJB+4FbDAMjM/QN925xh5XTjFn6MNb2q2yn29Q7L3rCuZPQrb4Vn
lEQirmTxGZ1E+vr3rJPjXwz6dreTQb/ZBO4iFjveuPzjMlqJPyzHguB1VpgxGTPN
IqMyha9gI2WVCxiYdOnU3qGdds73SXmLkRRdn+veAxtnq3kfDb9Dkm0Mba9yro3D
hqg+l7kOuLXNiFKheBoksg==
`pragma protect key_keyowner = "Siemens" , key_keyname = "SIEMENS-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Nfof9ZZHl85LF7VV8kwqITImnG3WEZ0P0YVzEeGvnS0PevbCKwpIf9HZIn40pDjp
6C7dsnYUSjkFk098OQT3cxa3sB4nEQ7tjghscEBIcr11fLIYDU+4+loBl7+vKhSE
JRtG25f4RN7VbiA9wVAQvgQi4ruRsPHC7WogI4wtvEQU35OHjmeDHS3L+Wnepjea
LnfRJMDlzCoG/Czx+a+eVXCSIDfoPGZ86v2+jnHyFeDiO0Vs+tyViM9ODIUyuDce
hi1T1CYfxnmsbjBWvmVUO1sVbRzXnMCK18kgayk/a+4zZuMsazRunqrSBabjCfrv
HMYPUZ4HGf4jWmz1yLuexA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4288 )
`pragma protect data_block
X97EA9rZmQyVSKGVAPf+pA8CK1o3C81qFxKfRs0qOQR2zH+ydX+N77GBC70b5jxR
f7gLzUE4q3PYwrjcJL7/afdvqh0Pp8v/SNilbMnD34mjydvwzGjQnDJWuka/jhPI
e5SADgvXe1boC3wo60+VEEbdvzgim3hjcA7hVhnxhD9adPktzNj0IbHZc6g6XEjk
hXbjsrqbLt9QQ9jTpFY0Sl2YQIUhmZIYbwdXZoIOAbx+Wo1WN1+7JrB8skeHjcBB
Zhp7ZxC6R4Ve9wLCBQ0Y1kXORFPBVAr3H+vA3NSfCUkNDxKTkwsWABvMmENIzfep
mxUjjhSKIBBAaOMFFzqczgu1TP62P2uqtbbmtVZc3IGUnNNm7gb8E5XDEMDK2tuM
4AWtjwUpVVik/i7gAOI3zFboS7l4Ang4YE9oimWH5Ag1IF8fkh8ebM8Gm+TqGoRV
W08t9OJ/kps369wuNrvE8wTvDmIkVWmd4pLEjSmrEjKDAcsK2dAwma+u+crNEang
Kkv1I0e8lbMp9YU+d5rjgEE3czA+69AZMW85A0WDYUtBNzVWY59ipJkXCLGt3/B2
m+5vFKdGvN9BdYF0tFZl9WIbdYfNfpWz/yLkzD9HZDVCMj1/4rC+Z7smZ3zAH4Iz
ejonoDqTaJdLJtvDaizMubBK56t1dfRaFNo1lOI13oBCnmi2ol/rYegDtxhJtDdJ
oYCHI1QUNhv7zPXOIvbNdJLs78g9N6ZxNd7MA/7u/3LkSyXUErR1srif3lOHjK+x
yNqmvxxQ7Wx4qw4vs5/L2DVtHsR9xNjLiBs+7sfPeF1E7lmEEMuzoifMdZztZjlR
vH/bDoaTW66nJcERzXcX0YzMX2vY1emTeSUzAoqcFDh89Z8kh2OJLssqkTctOWT8
mZxiZQvy2H5iyEAStPYAxYpCe3K3Q6ht0sleCnJ2d1aWK+5NCSaepAEzszlJ3P09
bUKklikIflTi+qm3X+Q4AONTsKoggFCRUXHM6uOIA1sunoMdQhL/pGcXvGovEMgh
R7dve5fUyEA00sQPmmO6lJ2eolbCMj5vHqJIefTF+gz678wUjpkJIwg5oZJwktRB
IvcsT+/vrSZCtCgjOZvfWvhSQPSSfdws/u48zZ5d8nfhoKxwTNWfzR0BlPVDyfQl
ekxne2nwD1UxEANWbbXjc+TwjAZws/QWd9stHGdzlE9RkS4B+8i+EibHfB8clN/A
jYtwsklGwOediy+mmKi0sq40l1ebb68WYSdVW6+ZfbMzBEij5e7Rbxbtu3M6sJOH
alqy+Fanh27H09T2xw3+vcmErU2F/FJS5qCaagg+OHaKhYgYIKhdwO8wF8R7L9t0
/74wl8MDZSvh07eXDkL3xaCqDPbtv9dAeaGdHvwnEKciDafXkdrboTAz7nPcR6LX
ip8VGFuAONSaTn8R+AZiG36ogZdhOL/KGPVHnx8FzwIJpYMxG2I4pC08giF1T7yO
nHMtA+JTjVQPnMCGZ0jkMICyVT+EI6wRsD53w4isYqve9jukUD9G4FmOR55AR9V8
z9b6iQoSoQcwlU1fzqanbFbMZ0f6Nqmud5N7xe2DLzIw0LxoGo2Mk60dZPNJQsQB
INQOdGVly5oSNgRQZzOVsJwqbQLTbkZtrIa8lv/PfXf0iPa6xnfpDbdwkNnt7Q+5
UFBDpPQXaKHKt/EiJz3B1uspdPe1xfAoxzUOgusx6Hkb0kd63lKC3N0jwETnMCUL
PBCHnDJGRZphGHTVE8ZqL5ixKhKi2nPdrKO4Zk5sCHEpR2eJUobipB9Pg+wI918s
Z2X4+XeaTmMyYbqUZW8Q0O391gL8QBlmI2bedJp0NwcgIjbenlc5qIs3CYlFo0QC
Pywv5rSXuXdDW4V9JPsgj+2zX8ciiM32d8zwloDodaOzBxp/et5Tkr7jMMNPA3Tl
6Tlz5iA8Zt4jQ+e+qc/KJzRmBa1gmCG7bymv5XIYtKKgKOgv1+byxIdLYCMZGhIG
7kq9ctIXUDco3wC8mG+xXBWE+osZIx2b6l7TteZa/Zk+r4XK1ikGo0ukN71wN5fx
E3W10XsFdVVV2fp2LneAJwUUniG7OTicH6VlEfMwJkFMEroA35BFiiTj8s/C53Ap
Mcw//CzsL22voXV46MhPjqWAlbWf9JB9RYgGhfFi8pVVI2tXmMrZbZntavcYCsrA
CnyteYSgnniIvfLGWAMi+y2KqusOLETAjbrZ8BdN3fioKcQEnR7Qe5ePQlLKD5VE
JusFOYxwc7uV5TAYk2UYAdJwY6MaMq7Btl4SYb+UsHJfMhTbwwHQ0zsIW2x46S4A
CfVI9WDX6PdzxPCnYA3JpiAGL1JIHMzBTi1/l5yCJrY0lzJRAtd/RJELxaDDLbkD
Yx4+l185g7ztYG84IFaxpqXvmSWDkD/5t9w4WIsB31I4FcOyTygmVE5vJUsi3u8N
nqfndnyJ9yPmcmIQobA0LJbgxXvJPQsfWUcL+kmzwtzK+FcaNPvQ8lkkar5zHKlz
5RCyd3TKySAnX4q5Zb9I8Lg7zfwClUA96Hx64uepwonXw3+fevJ27HMDyF4rEidg
VKKKsP3TYq6/a+6U/UgeJe9GYxqzCzt62S1kde1TprEdw431j8t/f0cvdMwhRwhQ
rkKWZdn3lgqAWTCLhDdBtIRRebDauNv92PclN8Y3Q3JRtCXF7pOJ2KBNG19oML59
i7z2LcMUi3JgWWZyiyOb0JGY0En1BZ197wJqVOPMesOMNc4AeD5IJBz3ZLORlzAz
Rq0By8iVOJ6Z62EeqhbBv2KyTj2P9q7IgQDN4pvV3pDP9vpNxVq9DW9IDKfTIEFk
n8g8tSXRWE60Z+va+09fdi6P1kh5+YFbqfp5FSqcw/o5T53GjPExWUTJBaRFsPnQ
6gF4Vrs92wNL5MmVED+ZzowDz1N2l+7mT1s29sLpfUnS5IE7A05FNubFXaZmIyCK
oJH2DXvC0QJjocHr0poe07Box1/6w8gKGstjDRjerdNwfnHusWaAvx4nZorl014+
uzfSsqu1qFpqiJbX+7fB0F3Lb4VsWNInLYVhdlpm5aXotLsTCT0KmnybcTMq4Vs2
DqZJz44VhuauSmbLT2Jq9FReUGwS+KKn4/JvLAYuHAO+DIyumkexkvFPT/pAfajk
o1DMEHsOZLjcid1mvhgGiU32xuW8wC2bf4xVuSHEURLf7UIK0jDX8T9BHA1xHdBB
fLtAEa+jVTc4QRfBZgFYp4sNBwrXsV9NAKHV8HXX/mjketCpFv+Gb6sqQb/FglxS
Yh9ApKF5n+VnRxqNAxjhoBIKRbxlc/5KQ7N6oD0APL3I9I6oocJ+RJSgEk9fpLWi
sSR+HS7ypXxXgxmA0gTbkgKIABNNwyhwVAF+HU9vohqANOEJNygP0rzVDJby4GVT
llaMRSBt/pmlhEQWbCxbdb6lWiLEZLqlz2T3+I0PZcytL9LMW3k7mHKOBSvsscH+
IJHl+0m0O9bfRFlLCTPBqlULLllnFBqyLL3/kbjWjPUwMXcnFT812Hd4d4TcVLZw
CgifH0Azmw5Ryr3UH6XXzxhKgQmClij2YA343z5bEDeeaX5JfyhieSuDxd6/dpC7
X7FxfPwWLX8+Epxwj+A3J4a7kuxIv8sTEkSxFSheaL7BQYQdIbCw3fFqt5gFIeMq
YhBGKo/HxhVrGQuyep5y0QkZmH0lOgEf7yv9bz0iqmyTzxO2MgeUiN3YCg/6o7DO
j8hTdftICEWV7jzRjeG6KPuj60MNySwH0qiKga/FVbHoCCgCnbCJCVHIJ3V6Tjli
ODasI7wvSBWfvOcVDvcQhtE5GfDS2175NHA4e5PS/R9nsRaChoQYJyuemqUEp75n
LvoEVvCuXx2hHeoiXGCJswKvi0Vg68bbl3H/VXKpkFfp8+eldgVjeKuASbynUICh
8qnv2SEq/JZ5NPsBxy95MAlhqCaAT90gn3xsHzOSaxa/D1FUDYANVKYwSGO9Kulz
XV06VXPx2G6YydPkmZUnn44BiFtQQE6sHTM79reOqOD+5/zImBk/qNaEvQVsVXfM
nttsF2vp+/HTHQ3CdM6PoLAdukOpzkDzNzuaj+mtHT6/6tfozYzvE8XV07UIQnG7
sW5kEH321LvAxuLxT0ItIdE/u/o5NRPUdIpt6BCW87wbOVY4FFuHrZmPfxvjR/cr
GY1wWkNjB697HkUILocXAKx8nJHB10keO1bRcM0yC1mFfssRdbrg1xLxrJoul2Yf
mkhiGQjApD7NAyYfIOzQgPwEDQH52h/VC1403QbDqYIUVlgycPg67P2qADS3ObbA
tDJYWCp9DJBF3Xs0vmetqFM67rxZGAUuhGMGRVcMpFmX7s1FVaVv/7Mr49POX9XK
mv9n9MK6S2rSErofHE/+9xsFLS43U5azSwTgPnMiPCWHeFc1SxQq2yJR9tqJPhPp
8i87HNvrD59PyT6VbT+5VZq51Bs7/t2gWDzFt+owA3oYYckdo3nN6bmYjxKKmHtp
mfmpkkYG2uLehgXvZT/gI5gF6sIRh8Mg5Otdcn8OyHTOq/Hn/ngbXEpbfX3qC8r9
S5XfDr20ZKfs6943PqhFEccWC6siCvFGs6lm6L4R3dYrXgXlz6Yb6MOgP30GHIYh
d5W0kT0MpAaXP+zkyz6DH4OIGCIwY5BdBVPhOfn/dOqhsnnmccZdfj6RVYXK+YIt
Rd4sQeaMgaAP4sBIk6sveA3wQMKv6bfJiH704yy5yZnpXw/ZZQOmSAkspV9fYYYQ
mv6Guobuxk+KdlDcQ+WK7jfKVgdAAhgbAyh5mtu3BxXMZ724Kf6WYwa4icQ7/83c
BUp44S+ljdSRYo7n4speThbeAlSlcGGMYoXaDPJcQHpzAVbcO+/JZu8Jwpews92x
wx44IY/hTBZZs1FL6eI1WoqxUH2IStzOLP7MgdkRIKdCUttNImaR2OyEV3CR37XW
zhRDrP4m3NMj2YxAvRqAyrmzpv/bfNmTIXbLWgeuCE2Nuo253KqMqaN0EBoVFs0T
QfivBCQhQFx5g83P7GZQROaQv6QzRfSyPfEd/OnsX9BufCjiOvTWEU4U1hsrr11S
pUrGDscFKXGQnlRkn9mhWp4eflCwDvdsy5k2E5EMV21opUS/wIybVQY5fQ7wp+as
8p1bLj5pC+pxDt+UVTbB1hKE261Hzzam5EeTcjb0A8jadAGZ9pycWUCNtF7UCBTX
Zaoz4bCQjroKB06VktHvDciBF29valOeuz08hVAls2ngSydrAcEBvXPwwwuKX9tR
bA5rRpM19xXDBUk5NEi8sh/vDyB8d3y3HcdQyEnlmOfDoloY5Z7h8oi3ilcJQcGJ
8cOzXarjODunJOVygKDyhZEca5EWEwDkx49TGcPAdE5Jnw39TL5cxac3ERxX6ojE
ZgR8kM6bBuzNVdcIQ/n6OpktOgcpoqb6R8Bz4iUb4zVBGFqkrYFGyzsbtVn9QtUa
jhSxj5FiynXJjlVsNNlL/1ZVA7mnXXoBX4cX2Fv8KDev6NLzqKPwYbiIz24eI9ya
1Z5TYyCuP/0EZLdPCNUZveNY4RspJFIQuhnOSIvPGDTJsS71I5beJCJ0bur01zDu
/Hzy41OwhFkW3GXBgwtgZqThTXp2t8BPdQfiRjZWFL/frfzCkCRdJkOY84Iyugm6
e+X3is4RzltxP3oHsgBfyBxTaMedsBhoQVW13478CX2kPGk3oQ+xUgfeKpwDH6mz
A1csd1tPOJMVvTV2UTAmlw==
`pragma protect end_protected
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
j0E37xRyiRtTYmMlyzU6UQV89YVbreD58sIFgxU8eS0jOCO1DACCMKyMmJZUvasu
qezU2kiYq8BbpZ4W/l3IKSSwgBdif76LDwPzdKnJH53WqfsCDwtPe4Sd/z1Nre1X
0b6gOHipbniMtnd6RnBzx0Ymk4Yg0Yt6n6WQnvq8O1z/qve8ySiBdREF6Hd/bm9L
+5vozVxzOdDJGYjP0T7bTGMqw7RtODWxo9mvv76M/FQbYQBN4unUX3Ti82/4J54N
gZxch5EUXC95/AwHOmSx0RIQfa7VRY+HNLDYgThnnc6ASfuLc8KjidymzBbpkvcO
WBmH+Z2n0KOzNs/xlKZa1g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 31328 )
`pragma protect data_block
vaDCFERBuUAKcA20H2VVkkPKauTRRKV+5qYw12XmwCw7Ni0JSfEin/awkZgQGOPt
ytHdYaGYr89IIg2KDAZ9HzVR2dSA3eaPxWTiZx5kpVZsR/FZI30U7Uik0AU/V1SA
Md3Nml0KBIulJQPESV/h/g95oZGPaO6jWeAb8T0EiZXeYbDMg1379J0rA6td+TCt
lFng3o5iPQ/RTKGHONCp9tuCRqLIuCUxtHPnPCU1qKQsVSXo//0jCTD2Vaq9Nct0
pMWOtAEGHPU2c+XwofxQO4VXe+shwIJ4GDxAq5hQnw4imXH9chVwtY+cb4b7I0Hs
T8GunzHv6KThXJZiybR4gJfly5NwMkmU/fGLMslMRjxDlYLD5L0PJgZ6hn7qSiD0
1jB5lwnrugb48RweZ4Ne7Can8CRrdJTlYf2Md0Gje0s9IPAWYUE6BYrHglil+89Y
g6xcqk8ThNiVsqXAyRFXFPwt8j15PwUb7D5UQExE9vkiXfPPbIuVzzc62AeXtzMP
uYZiKisfKfR6wQGZgxm8Gm/EHlNQFKT68WJrCY1Pz72kaTW7WM1T1thsneXZlLnH
PwHLwtAFOp9O0Rl0x86JlJDqLz5/dDqS1rUW5g+k6p2O7bGDl9HjGTTDgz1BtR8L
WtK5AIByD22p4/WDDnMhEC2z0/hTA9+a4w88R9DrcvpFAOpHls0SukKIBdiIl3E1
GAkYQUXC2xAVbmKXNuNNYQafti3a8buZUTKd67c+mcAns82lqU+QxxHS/bE7EUxP
OGeCKIFdNfLSG35NiOIt+JzWXbxxq5oammuGcAZs4DamxtaoI+KVjTI8A7SVLgLZ
uL3939lBtpP6Gf8GCH2QdwKHFyqvuuemTTmewRYD6AYuLJgWtyLyph4Apvg0i1dM
GBZpMP6c//ZmvmIgwYZzy6fvkoxnopzuDmfz9RbuHJAKZ6tZcH0HxzD2eagfBJOK
AK27XK243oIaExcuRcCdn826Fv2hstl3iNioqdHzWDYjcqcr5prgUPmCNzZo7Kro
9c6JvRpZubvAeBEZUdQFqSa+RkiSZqUmIfZzfdrXLmK3rqwvqnRp+B665oLWfUEA
DnhzKE0cen2AuFiy9BcqiKsP/upF4KoN/JCbOJoupFvm7+cHvBnJ3xuG7ASAKxzZ
oJZxKXYV7TAvcRwR4hROSAWfKCcDtVVgzGxc+PygFECVDkHK4w2OaHXqeVNolbDG
1RwDo6DTRwb6DJ/KnlL4KLIlEqYVYfyv2YQ7wNAN5muVwNeXkuq32bAgIk0CwqkJ
sxahrpOo0XcptjbhRdyyMrmyzlUfR3YpC2aAc19v0jXBYBvgeFGUoX7iVMb8oq9k
DSmgn/YPNYimo9rJBRQIKhelMNfX7ZcMMyoruFzO9BFyM5bmHGAOfe1Zrs0RPuwS
jSYWji3tosqdAkCFKsdutzJ8F0dn+rYQA1HoGza6Hsqb/GS+6sdtGY6vb5h12Ati
nIHgibl3cSaW57ZXq8SKsWfZ276CWpb1Rs/YiXPL0ic0MLuSTjK3p87yQ1Yrm0K7
k0qagBCPJNpgxujloX7fJqEr9NXfW7DBmmpNDDt8leBdUdhaEUvmO4HKtffCzOUo
pp6FcSUNH6wSXC++VSXfP8mcFOlBDfUmpr7omJRF7ru0+C+jRHKsbEfoAkm65y1X
qa+0ieww2jDpl8VoIJsACWTjylfi1gCY5Fap2amP8xXtIVD/sSijBCpx606omILb
q6rzmF7TSChJx9pAKyETBQhlQckzCvptbxz7pD/ICxkgUAaR3JqNfVDx95kLcW0O
L5LY006Kf/yGZTOc7qGZ0vE0+AdncXVzVSmJflziiLitrjeA5oksRSiX59K7+l7f
7D4yrx5GoQ1flEtK9QEQJ9bX5GUVl+urVNLTLkAw2h3/Wd4cpOwOY0EkSie7reae
wbVwpmOCskqxYpWo35/yoU1tSxY7iiYRrEjvKW2a0SPBxLFnHkyWBq40Q76IwjhY
TPpxsOLcYm6PjNRkLEbLmJVmP4aWaCOBy7nz9zeLPoIJULkaPNTgwkygrAqN8aos
STd90NX7hF69laPjH7myGvOmPySq63snTN+N8X+TME75Z7IBCp4EUZvYK0LghsQj
QfT+fumkzCbO4Py4tZd3WbujHXkrANhQHAPSKujaOrVO6fAH8RZyZPCGS0UVMXDi
/auPCK9xxi0uyvenRR8z2NLlm0lljoEwKS65HP5e0oKqNy4Nt43Se+jOVzAxfTdF
MgJJEXaWP/dHzUU0NbYd81gytmWwcE3kfLO07DJTMTQQ1up4RpDI8JjxzAa1H12/
dnPfEgVu+4CUejizAal8UhcvF/WEs4sBq+A+DMZhxoudICm2yg5sF7MN2x4qy3Xo
QMa9UGqfQCbuY2VPwQr4IuddA0Cg0yur6ixPhPItO1BlAXLgtcfcUEpyBG3dWKXt
wJrLV+Kopv1iAa8XMNCcIfcBjN3YmWAlU6M4Go8qrEmMIZ0jwpReHX7GY/wP+iAk
VnHZIMOtyD7/juf+xL7Thv8eeUiHT7iO9TV4OsEXKTl3c6pJlkJYOZH1f+g0LfVh
lS+hkez3U1SYPcigvRgx3PLjVwlF1nGmwRkLus7eRd71s9bPLjY8bUs/IpYHtKG9
5mMobVw91rLhPR9zPMSjHNs7R7PNpXUajf4kv23TZhm8mGHkkISYrVPApsbRKnEX
A+NwEtsRj1v81qWFtGc14yTxciaqhd/MUOGUm9yDixX2ZTitprq+1adOxiMh2uR1
tpGYOP2qAq26glvoz50z8jnp1IiCqhK+3/bpHfpWdUdt9qDRyW9UnGqahssYBJxX
5UfSAF3y64S5Bqyf/0oQAt5ukxc5gLduGuLanFF3C/s0wrDaoQ2ob81ysR24k8BB
D7sZmjOmdLAxv91+iWhAuo/mxI5HQT+ZMJxX7fPHTmFjgtwb7Sv6aQ3Pl8GBAi+x
vd6Axkjxe2Sky+EHl3J8UGiIuc0/vNOl6fg86aGSqrFxh62d4/UAPZuE919W+XbR
ksOQq/snxlDpyVcC4r/uG7IVpiExOxKWh99YSo2mOQw9yolMYeaGdVHDN0NxXjZF
BfBQEr5E18QTXRyOZlO3edRTQYNJsER1c/AQvrLa4v948tvuHEE1H9c4+DEWnXeT
hjr93f6fuMgvsYWx2laGAEQIVTVLM6+2DOyFbClKANOy7ZjyB02JZvPISV5Kq5KS
akKTB3wjktii9uANYaW3OL0gjE5InLYfDgWWcDhy01WFZJ0Ym9ele76qqkanuE5c
famylnMtikcQSqfcUsskLjDZqyPo2IxlxZAWeN+/al/v6GfNA11JFJ3Jip6D9FYO
gn1WgUANnyOC52v1+SWHS8mA/NSLrzDorqB5opGOCY3p1kIpKx086HAPuEpA9+IQ
20hAuXpJOKU0H1Rn9P/IGZuWrcHm4cEUR+H14btLioVVYZEZRjYq0DL5Ee0zdjEH
bj+boT1Cd/xp+ZJUAtUYLM337NvLoVYoRj+r55E5/osQJzqwowFc9y9zywmHjkYZ
eykwFxVKIC2PiWL10wS5mV4vPVbC0fmbvI6jrJkMTu33ecRq2qrAbNvImaouG0gf
2iZV/9ftbDYupHxFXsm8GtS6FpReHRgtlbLWZsN5nS6YZ1ZQaviJdKqn6RPFbsHQ
M1+tqG+HUaBGzNawBA8E8WPJFDAorw/Otq9YvcCAyMxovWzWOuRwVzYajd/zvy0D
6mnrmdqj0ZSintvhcOYZDDhM4eYQB0nh62XxRUYjpLiOlEuYYk8I573u5W1Kv3+6
uWHK3rtEcLPcySbZaGK4UE51tL64a+2vlFeNNgr9Zct0+IcwXHSSBtn4q09KzIDc
1NPNq2lTjc2xERFC5b//W/xCTEAazsXDiN8XfZ0zsoeJbX7BVWVlRZ6ryi/ZrRq7
JqAtTNJGN0B4nWgHWh/VGO/l9Be8LJzDvxUfKu1pFgzHyHPF/NMlTqcXBNUimvRI
eI+2N6nD93Vbtooknepp82y2IFG8n5IslJnsQIGuav45R0VaZOHE4B6KTauxrgGE
RaG31IRQQ4H7nd289WkqX1WhzeX8VxLxBuAOY4WHk4mW042mIsH8z5Yw+34BB8s1
Q51/LJy01D4qzlx9WHw8gZonB2bn4B6JxSPXfB3o3PKbst7y6mYYu8wysd22xJH2
VEHTgvYcZcqvpnZZl6jvjtaY9yb1yRpd4lHWIyslWRVsvS2fJtbZMFl/8nPhCkF6
UDB4xvTCloYEHKXoLt7t9tAyUMowSfhyHYFX2QLQCtYMAeObc1gSP/Gsun9UrF/d
PezeUAdIhLNOU/2wjY52WHwfGx9JGSBlFlQK5A/KE+pQjye9DF1GQ/Lw10EAquiy
hgPdbT7m+pm/wd2HFiHRfxR6gek2inAnUQ8/OBPeoB/w0nE1aCn6fyvbqeBeggWY
XT1VgLKgeMQSsNcALF+HhVbPT6yNTDKb4bvPb5Jq4ROIzU5qxlwwMZflS44M/Mw/
22I3SvBHMhQ/9n3CH4Jxp73EAFK3yFZT8Aka3/wfTc21E58idzEK7MbCIpZJjm9x
vhFX8onptIW9hIxA2tqj59O0KDK4pc92Ygf+aBo/c/xtb3RpuHSB72jhjc4vZxWp
33FRqVmI55lxPv+Uf+stJm8p0DW0CDcnSJ1KzdE3tGl1XlBWuLE69qt3amnkjgSB
NDAV+uowHMGot73rRre/YsFiLrfSPaUuxGrtUfaxM0TLX9ixmK6qXCfqa3WwpErE
FiFKw2PEpkBCAP0+chRqY2Q/q4vK9Ch1HLQNMLl3YS6ha3wZcJloDPNOxxLEaihj
5Ndc9GOCA11nsGGfmctnaz49U0NWwi1eDQI0Q1ucYVHFb8llUFhB+mPK58UAPZg+
aUrqzeJWQvWS9FuwiGJgPA/7BiMiA6QUruiBY4SdkEq00twAihtHv1gsJi4S4gow
6HHq+l/DLW+xX/LcQMCxRBZLFVxSFZLVsZqkoCAVf1Xi/IB0gBm6VxqG76IbKCbe
KlD0x4uyJ59efe8BLolis1SF92j5wIrZUTaVhOHVuGE7hXbFxxC9TOeU6RiC6Pd5
6eL3GvninA5wsYnJ9bhH6FK/XXUpBBLFk4Ya1TY/OvcRhE4bv1l4c4ECO4WpeRFV
fCgcxURPuQs+H26onthTCmE14aphWz8kMpsyyAxURF3OWzdOX8aKdIE6qKCk9air
emSyL8qHMjhdzANdIFp0BDXtgnNYXiDfRv6ik+4scL6qSuq6ZQJ1KXxg9LmcqJ/i
rztAvL15sy1DaDOw89gEYjlTYsVCR56ZdR+6sVz/v6qBrZUN2ivMrBxsYXDoOkbq
iN4QKf6HUPS5VTS3UM5y9WeoLJSQe7JAiKp6lLbphRFDiakz45j552W42Bmx+4vG
OcvpImqdlJwOasf9OHE6grGtXlAUU8ysJ/D19fHx5MdhPico8j27WKEyrpz0+woL
b8ARlQv4hJAe6p9wUVXUZs15s7Bv/lOJ90wEhJelCs1o0JFSeILdH1HfdMrBEEi6
hVzhDj+PpBuGw+LoaU1yYgamo9cWFXC8eHQnbDo3ZzbJqnv7Bcyfc91DbQJWslBt
as2/svvKfda9hrkPJess232r5vcDt4G7Idb85OUtj6pq7jgvCCqwRqiDP1Lj91IM
4bcWB/bkBEmXn7kdwnx2fYfKTiC2XMgG9fta/BmnQCHESu/nqw+PuJpmPTUPd9RQ
w4yuqHycPgpZHlhx9Bl5Zr3QJMtzJJkuZLMW63rGmO6LM2vhUgaO2jUI07Jan4ty
zygPjxadmwmiBq6kEYuzzrUJ3q1IOHgDZH0JHo8NMAH4xW+CutON7KxJdLAmMZAU
aJMm/zoFoh85orMoN9qDPs/u3tkmktoaZSo/VH/9s9Vn5AVFKQRKM8yON271tzsM
Ee3vrnwunz6oSeeIKUs1SH9pAvJx8WspFhyAVBiyYXlrGIMT2/hxlR3Xo22mvQjW
SC4xr/bFxfuAISx23Pd3hnx/DpINS/KZx2cR+us+RYC6AIwCQepxCwOPmY6n4VRu
/gF3I9b4ERVp7NJ6vIm9J33tlxLaW7qDSyV+svWwnGwy1jUeaV7YZs7ZJOt07Sxk
1ZCi8Ey8BpzcR1AZEyIsUHoNygYTMlpFyoDYsX/wGsX9SJzOzj5rPtpctjY4xIMA
xLsySP98zQOqy6T+9GJpLvjPqUwhV8m9c2idWR7SCsl2rJm4xLvOwIsawGVAVU6I
yoyxb793QbIT+6COC53Juuqi+wRoZXuVsk8R9vdeT2/8N5ibGuERFpKHpW0SSMYg
eIRDZkTZWRxP5u45d1hh9CTTrHTRxlv4tUDOvMOv6RqefOArKze/upe+D+Gx1MtD
tXLUs14tZqhbFEh9VmcznDEU4ydbJoRWH4NoiSsSqgitXrDaXDKHeMAkkdbfuAIQ
EuLpdCihb1pZas/mEuiiPj9Aw6hR3C0SH1KyaFsCmuQqlTYnU0krxa9iilUk+ZIA
b+k1kCu5lm78wnWnjjAFKHB1Nqp7a5GahRgy7xUGeCGKC0rEZhlRKn4d811ae8/k
oJFPQJjT5mrOr5vhe1Azrf2M1ZJO8+7JA5Y5qaXfKwTlfEEc+cLTugrqSaNxF6X+
b5IZqCabe8ZCnrE5/CsNbXxngnYiHCjXsgFlfk8D0bx3sy+muNbfVLFyCvhYlWNG
zGEVdT45QHw5I+RUfEgsYdUSX4kHAMK4R6VjKXRKaBpEZhQeopyadDaxmLlnwSv+
ae0Efeq+vCDbgVSxk7hsRowFOuZv6dDBuwl3eFQ6Qm4iqgUSqyOaDKbw571ICKeH
9B/iW3Dhv0M9a4NNq8D6RUHtH8yeGn/v1x63q7CjrCVnLbm+XgfAgxVmzOXbGhPj
jOSoUAD2yfMEric79Y5XuPwQ5SYtMC429sIj0U8PocFdnvCQuh7KwxSqmlGRKsjb
364ogjxHRb+bS10XxZfdWx7tvyaFk0q5ZX6yViG6xkBuwQbi1GUf7Y9zKq/6yVH9
aUmvJqjjKphFZSx6NW3uIrH4tpHl4mQuCREjaaJZS2kpXZ28flwCT4beDeBHoZDU
1bnHkgVsYFZTLTnv9MaZe1anfsyi8Ygj23be8S8xVuyPPuUX+SFa5N2mCpJZVrgI
1sT3Ky1b13leqR6lqjIbPo6FWAMxKpafQEsiSmENlFeEZbzZU0j0Aq97sbe11MMu
/SQLFkJYS+4CjDn4+QTjYVB3F5G2+ZJcoeBA+UD+ovxyc8eOyOohpheits1qXGhd
HtTEEtpmom2/WzkV1RqJ7CR4Cj3+/1tk04t/xMugGICxN5qwbhUvK+7UwshLe82X
3uIwrtK1k3Q+v7ZORVYEBrIMw3PcetoJM9+mmZQeAMj3Alc1Ws6hYgdW2g/6JOvM
WlZxlCmvjTt/P6jxt7Vg9f3JOB2um5wmhKVHuG2Mcna2sgBqWB9kqjMxGrerl5gS
PO4CR4Ts6lHT13cSuadNlTS6n/izjsz88sV50JAhkWNDyB4LaxnISv+YjK0wFD1k
w+ZmSbGslWLm3Y7rAbUvhOBjG0fZJIOSlpOXYCwdvV3EZGxYD876K8GW2Kc8it+O
8g6MYJHJVUfz6TjfUr11lHsL/WYp4dNWBXkhH0WiqR/QgLRA3Xrzp8pEGne8pf2h
lSBBwb3cI8LK0I5khGrRXx3jkDWEYcm/YlR2xpdRIQ7opntZ7nz+I+PTht7Sz+JC
tg5i3GMvn7UwKMUJFBwN5HGsDOBCcT6tMLFNZ0X/5S/+Gtpugcn4kXIk70G4vCJm
pWjg5X3cM2wp+y8waaw6drSYtjsLV7osG+Kd1zW9Ube6J9TCGIzqBGAc+6TU3mZ8
hM3LKDOc2az1clUHy9uZV9Y1VbK8gGVfifnrxqlHGyktrIPaFdE1rAFCgkCpgaBU
z2bmcttW4KNso4QrlmUpXDu8GEmFL9fQMAFaSAEnmMLtS0SiSC7HBqwyVAlxXhMZ
+8GsBebpSTg0HCQ1ygqHUbTPQurDon7NdIkHK37LkxXwhn/gGoNFw2N5x7KRS2z2
vTIjXnzFEP8UKAjdCDUbKgjKNObPjJUN4JV2q7JCASaHPz+Hf2R3Te39h6lwWkFg
MH45z2ZT5m3kWRkKLgRPLY7mU7ZFv/vdMXV2F3pFRTlvKcrDLMdh9SGyqrRLRcdi
ycAM1uvwqdMuwzCZrl6wtCe6EsLry9HTmu40S56EnCyhJkgMgqc4qQafCiN3KHrS
KaZ7tr42G/RwoSWYLFkOtelFKjvA75IWFIghr3w9RaI8qNOGQUq5BaQkg6h+EsHy
NDQIL7fOS/+xq3/1Gf/k/orCU9o2WgGkTiyF6m5eYNMPWRa7HiuYPoyeJjfdW5Bv
Xc5F2W9Y+hmBlJBVSZGe/3lVFcsEPIvvN4AqGu5dPXHqljaTaAwQR5TuvlWzOcal
anKT2sfVNb0cKhYx8rVGpszJ0Dz6RB60PPrMVbrTwZY5MPZ5uXni7m3NxnnDmKUG
G9p8nGRVNUuj4y5M7/RyDnPswCb+zxXc5OeBlSNA1O5n7eD8xXIhh48+oxvRWcwh
SbTpqtjN2wPtQEhn7YitbfBLplJftVWq6o/xCReiOh1Ig1l7GQW1kAVkF7ACcZnM
NlrUOOvJXiGxaIiTUEceF236CUepv3S5AUTvDyY0Bu1wDZMZVGhkiVBiNyGCYcHy
Zo8ogRpXrN+rGPsMGGCTPpqwGzecq1vmOwJFp2f6qpesSQ4wD2Y9SVqBjxnmFmO8
Nv1KLIZDsvcmEKMzFfgqtTNqPTOZ491DzEmMchMthYu2nS7gMdiwIyuV3nAx/3uI
I63LHeG1KaZsUNoEcNz1k5BCcUypwFtt2/FSUYqIXZdS3wcLID9lkvDgaOMkp/lF
dnCG/Txeyf9+ctCrnkIIJxy/1pJQcUHJi/MxBmhqYlFTpNt+1KSWuKzNTC89Sf7s
dFd8Av8smTwjqMB1mLfzmO9eRNPUIlAsr/ha5YU2ANLSeC3FjfikRWLwfnDGQ64i
2ytcAcdmMBPlTtkxskZ93ogZEBfq4IbY7oNjZM2OVNSYFdtCA/WvDV97Iy74w4z2
vduiXQWPVc8Kd4YHSFdxoz0wtBgXO8pjasyTfNTPo4yessQY/JGuI/afMHZnmzW+
nLmTFs6vXb6DJrIBBse11uYmPcDs1W1UY9Ss2WFN8AvLNJZdZdGGfumKeMg+rHHn
fF2zdlR2YZCPDT8eMw4rpBsNgoc3UW1ygd39xoBjxjAdWzkC0mW0a5pEhmhCCuPC
8XlqpKW4M0krJMfnVpiH8eW0eZH9TUmNgxPj6zDwnX/VPgLAOYwpH8Gl6ryAlf8f
CjK6dr/VLjCF/bkm4VUogSicK+JCZvblEcJz8O9F4KD1Pqh09Dl5E/uZdoEmhU7Z
PMixOcu4/V88QYuVqoHv5/hnp0eOhS1LhYKDUgq4A9RZUJwYwJShkluMgIegqvW9
3uFWEYXchhNgZ3Jjh9lA4lzeq6VDYU+h0uItXNb1w9krT5mes4e/otBPjrFMmuPf
KycZG/4eZk1txeBB3nzpSrHsIvmhtfDvQWlfu01whAf3Zl/EUEiHT/w6ogMVcRtE
UeyZ9pqBQNMdnhS4kstUdMyLMFpmqyofcPKR+heCYYL8LTJGGlxl6WNElWYdpztU
LjpbkD4JT/QtFoLNxm7mAONP4QmiFOH2AxZGC0XSWcRaGaYjPnS+tYBzPAD2qOPY
cZbwet8aJLGYucZRg5CIc+Ctt8Immk34WktNywzqaNwVc5NYwyaaKYtPM3zvPF1f
GDtWtlVgXYS7ClZe/EqNAKnfCASYIAxAylSdxfXROvjAObBXbdhGfViKqnnX6PrT
hNnrEqtBWF7dY5HfkZAC1VRLvGwJn9ZkF206AcYIixADTMbTrHFUGnMValIGOged
RNsqjobgAeTSUNB8I7flDCnsxvLJ19gHdttj3teIvFQb1yEzQcwXe0bC8TmwqPeT
Fb3cawYLj+rQ51yaBx6jEdDIF9TxZopq/WvGx7cEVo2K+zSA4DOB1/+yP5BuMyHn
1E2Bk1TRRleL1E4nG7BqSCFPuXEL5KOU0r6nCRdUOVP8pWJo2DcIrqRTtyl/786T
ob5xTxtdens5ecF1Ms4aV5DcLF/qBlA3E0IrzQfLCMtxSJQZXlNYHYfdLNfAUkAb
ipXpWAgyBuMnn8hBch69/+vkVcQ4ogVyQCGqSbb+Toxlkxpb9iO3BuqVzOL0jvAY
pM13XrAYMSEnHcj2iARe4GUt+BezM+dOp9OSmVqRcDSF00Srt1VGyAgNZf299w94
qQ2WmMXlN7UpGYWxNZ9/rPTWdWyzaDG7+/ybzOebRWCc3Zy02kaq4i98cpfUS/DI
JCSAsEdlvf+MGWqIrzrGhS+2l4HyprkhZqGgUfaeUO/qgB/9c1TY4mHTa87wcQoy
ZV9orU81LpzOFysJeiZpc/MggQil39jAneiIKE3gn1IMDlebCmXsdsVyVJms9v3I
JRj9GK0+PpL4DPClGsuk7CL6vEpjTPWGSTyb1q/IsF7NZ4JNW/MQu8Ir1rd6Xd8q
Ayw4ToNJM0fPc5bkgESQjgZzI3y/jIZN2FaMr4Qo5I8uaqi1ERuW0u9q7VV0cVq8
tMQJZREhJIbUvoTiELKc9G1mpf6L7abEdUKhng/Lh0fxLe/cEMk1zzoTH7V+xRcN
/AY1kY/GcbRFevPJ1F7fZsDq9PxmBUJgiyKRze9OwiFXe4yaI8lTN9MI7WoYJJpt
d4r/sXGEVeO0b3+1tq8yTO+/IA31xBCKkAdZjNLk9DiHyWOpYfsvGO1txp9EvA8O
+o5ZXpaEbSUm5BnEy8wqjPha7vNi+0os04BK6vrFM+lobevjt3rl+U1GN0i4vppk
dWsij2M/6Gt9eyPHLGBUMaBoubvXjNpIArd8PeRJoupdlM9RuaxJXuWwURgKrGBc
KcIf3znRHVb02ie1YUpnDvD4K7YGqCkyk4KMkvD7Xm2H9YbbkbTjuMXmuBPkNtXc
fkxNxJzVNirnwqhv3j1GGFozDYKr4XdGRuRofn9zSLObKL7n3Tz3iEMVH9vAtLqO
X7cc4RlRnoe7le5PK44jJV79cnPYiP5pPqwfaHDdVNd6XBPFdPSRsdmoLmbDAddV
9r1KDAf4NkNzYMGnJa9k4StkkqZZxpQFtHmd6Qm8JDwzhiTrlI6bbbgCYg0pRXMS
OJ5Rotj4Mu9Yopb/7ViE2LS/VY7gp3Uax1f0vMNC8Ku9LtCCc9zSWhP4QmEPTUux
/lTR89OYWFjn5A9nxY1P6D3U7UGHW6FngGyeoczMzlvxIaLZ8d5UNFHG07qNp1B5
8EgxeOtO6t8MxIANsNuFf1Ahxr8mRzbR87RjNs3f4y9DJnL7HVbUXdmR4zabyUrv
i60beZ62rcci990LUYY8R0tKCHLID3UWekQJP+0GyUE7gxoEEJOw2+2RB+PZ00to
NFNcSyDN5AQn5VMmDFU/9BYr7kUQQkFuWvqD8xHZC7DymrK+Utwaf2ErRdLfgTzl
YA9giGne4B5Oiwj4x9VmgCfHqe+2NmlOCJCbWzgDabh75+BYd17LlGtgUMXS0fJt
94IsSyfrGzJARcKBD8YtEPpmKFJyIoFECTepgCYb9BzHyogklKHM0I4ZOjLQnj9a
wDz/oWk4gogUrlFlGfVjJ9yo9bzRzoLADQ+hZkOAy0BkvWOzWPrmmSsKh7WEJH8T
n3rpXY21I3XkCUUtBKEwPvLzm9/KqGmfoOyn5hjcV0l/Cu6Gbfs86vHR0ZonT8fF
AKDfr+9ysmi6W22SKoy2LD68jdAZmfGJhrTzsi5+r0MEYCeCPW+bzkLyeqVv4Mul
L0swF00eKq2VjKWh/25owm8HeudisV+A6P8WeDTC0CwASqLZw1wfIS8mpssAKoQm
uAVbSNSgCEmQynrmciR+z0WcDcM3Ln3DbxespaemxEPHZTbFrsNzFUcz0+M6FNyb
L3YAEg9Ti39MaVeacd4gCeeEmGQW5VhQHv9pSjHlB6LgvqHcuZTbn2GI8y/Jw/T8
JcCh4kWnoXe2NyOVAROypeQIKMxVy7YBGh97FnEM2KMNeTAwEzH3rdal70GsLj+a
/BBTyPv340i4i3Be/dO8n8Q3QxLd/hWbXqVKvj5Nns0D/E+3K6WdzkfCGe+4Wc4L
SjY+zvZ3Ljp5WnkYuBPf9Hn7TnOHMxceaDC9+KuHiRDERT8DQ8vRuCzkC2azDee1
3Z3bHN2NVEhD9uF0/zRqpYQA6njqlcr3DFJ2Keei+rgj6NgifYufHJD1S675NZom
6sa7oNvjM0MgLP2qszv4rOBk9y+5TpHfUIumGv67AUhQIgVkzLbmSxlRYebAaQ3R
fAviWZl0b1MSDsLIIweHuGqHPuJ6hGEfMmOx28kDZ5jzdSRzyKEbjs5cm05YTVPa
MNWrc0t/JNldTRQtwTJzFU7V8/YDIKBY5RoFzn2mo3e8cqBHgbrVXExXQtpr11J+
IBmoMJ0PfG8E9hwIOSihmJQ5H4Nq9xJNYl7A1VZQu9zrqXBPmz72nx4hA03cmA6G
BbDwHDHUwXLGz6l4m8Y3Sp6qsZYIH+6w+sONBpWefheicxE2+4PKCppwCIex1Co4
aLWxGe94h9fORrApOCEm7S+gk3XL6ey5n8v8xkkEfqOeh4L+y+BLpDaBDDxHnivk
+MSHFEfb68pl0UGvECHKmRwyuEdF1NUIGXT9Cei0bigs3qpMWtvbChgHygnRn3G2
V1iJypqCVdClVjli55y1ZNMYF8DVOEp3P8U+tcf3b2JZIMSiakkrZ7XCAs3ehxqV
BnLgvkC14McbkxHez8YC3vqNbb87U6cyyl20ImwyId4YVMDLXQBH+k08sa2gndB6
QfEZ/+EMg3xl5UxWmvrcp0AM/QTWXYTfEUAjynJUQREh0wJ4cNYbParbjWaQ++B5
fF2LsnBw+KCalIChDb5oEy7sBrnLMpo/oeFn1b76DL3h20t25q3jcdVXGNdDIH5i
uqTMAxQq+4omcjg+rzqikZrOZEWMzGVnz2hkSUpsPlyFSsdvDBVWJPn5QiCVGYJJ
5m3GOceFOZxfGFuU1VPSEuha0zatUUCYpSXQ+Hp7DtcluUfH8qgidXmockFP0suo
wwjHOTgLJSdu3qWUHf5+bA0YQhfa/bUQO3Il9U9T4lfdMaEAwAEtzfmCm0SCsbrN
4QUu2HHfkk8Zz0AG0kyYVHYQCdso/oj7kjrk6VCsHiQ+82xYCjc6JtslKKmOdUoj
ksz3PE14JvSDd7RGi92vETRfloMYKP2sXBsLEU/tMJOM5osJgINfpTm0zGAdhS5B
HOx1Q8UOBfsCdgjBo2zpl3BqbYJpFRV9JfW2BUrgKlM58cHXEeVCG5+8wgysxWAx
7NrU2Z+8VdfWBaUfHofqWMFqUkregcnDHQi4Lsk2Kb2XbhoXHno+MgzG9H25iBTN
GyTaQVylq42F0r3Z+j2CvLip+yBj/ngY6aGxzb9a31aMmfoWu+ISncCZfv3UnHET
0Sh0caBsBvVectOK9z7pJU5AeIzwPNMcTgLNhHkFDkx3XCchtJWmbuYGLJnnFtE6
Kw9Svuw78OM5T67IeO28z103yBA3EQIa5tMb2Aa0hjpifTmrWjv+EZZ3fHRtvg7T
4wWTiIebtBZ1xJfFthNjWXGnuwEPU/eUIZ1D2SJNmVS2INkPlh5eGYg3Y3pqeIEJ
8AolVFbPy3MtLEmoIhaTbmMhzdp1q/x0ZSSnJU8We2H0Ak7PGtuLUV5ll4udBPDR
oCkP8BMI/zRAdw8WODCQAi352bNxAbdkvj4OJy8YuN49qQhTdIdhx1c+hnYrBJX1
85KcTxKdChuRZakRL0cjt4eB1yiAVBIf7XjHfGhnD4vLXAE9caBtwYHA9cheLYdC
fcbdkD6bKikp55JkeyMsuK3e3erRKsrMXCT5tiNChXWKuoq7PmBcjerMwvM68HSX
cYpQWJQ6q8Qp17dzDVyfIPQoCK3QhdEaL0+PLVl83La2iqurmNx4tswgahYHWIRE
VeZ6TwmMiEjjrsQZvlsZ0tuaHkY/zoongF9TA+fmwyoxK9ZBty3FKeBdOH5GQvba
ZyJqwVQwAgzJEVwKydzkK7wXPCHCLWRmCymBjoXvrYeF/zVt3HyYg+N6vP0fY9RY
zBBvESly6fCv7HBkahWu+zfNSKw0eeXowVFjtsQm3F3zk1U/138B9enJKY347zFG
Fj796ErXR+o8MWCJZaDS4EuNk0fh+QqkYRhNw3tI5PEXv3mVuvQ7i6VTKCYznqCf
QSfaTCzU+M6GV/olJwaOp7TJb8KCRyZEz+oqIyz1SseCxONfjONLI8+QXTdKDTgl
QO3o51QT/6zeIkgSO4l6DfQmEtNmwjG8i2a+Sjp+x4XbLMV2oQ1Xi57IAETY/hmz
u/lRLesIi9cNgAnzHx6exFoKWrqQA0AIzsqeVOBmKp902Nh/DG+OEbrd4YfjOYAA
vaU5daLidTrx2Nkw+egCjwzCsgd9EQYvlFBhcKi6HugPjmNVvfOhG2yB9e/ZARov
fjJvJGxRHZjILC9lFceiSeLOU0bDmqfiN6+3iKyD2kebagO4rCXy+nutbd/c7upe
L+5EE212z73KZn8cmlmGwLj+QB0Z1UERyCA/gqJt5esuivkJJCGePD39aZR8OFRA
scXL1oGvEm2Wq8YzTcBlorxpIBPPmmBvPXoW5zIjdMPlMRdo4hxyatOi663JHLDN
dngx3B1f422QLUtp9jwm0LAwbwlGn/IWbJC1BFRwAto4gQsJD+SEbfj4V2tcvpUW
QDGGEEh4S3haQqniPlfrOz/bG2jfRVehsmE4t6YjsAdNnR5UHXvQklrIKC6xOYD1
UJKtRju3lXt0tFWMnGh9S883l8qH/IKhb+6k0kMACmVGIdSsbKKgLshqYhbFzqE/
23UL6d+O4pPDk6D98osDBq9uS4EdPEwgkZZRTKD+U+9JfhjnKzwYt9cwlU8DPlbM
W9mPGNagnTeCe5TX6RTG9ZGSjamyywpIcgstHLaGPJKLHvJav7qLbTLanxO8pcXz
M6KzqJ6yFPvCht972Hp2MyTzXqLYbL7dfwGyrvr2yawGUQaBgtM/Xh3UaFi75TyD
qspeURFWSOZPKxuYf4Q2BnYwYdHUooFPjQT2FQpciPt/Dweq3DqzlSSRuHAwy4ib
FmCvyYsC8yQZ6URGSykC476plasBd+O0QperOzvGV/RcFZS3hbazsXqnThdmPngg
V4sXET8nAXbrUlcaY3kVYPxY9vhHuTN3lMwH9ngHIkz/cPPiTzxcMq0Rj5CUa5uY
ZifLTyW7p5SxNJk0iYTxuUxXySBIAlau3bEbe45MTKcIHsTOSmZPTAkhDP48sIIc
Qt8KHD6PEN26dXIFZxfUeBlOCSTqROBu9Py+rpcJIF4HFloxtK9SYtlS/3aLEF+R
LvkXnn7Z2/rkKmvNi4F1MwKzVGEsO7ba59dulDfp+7RJhcZwg/Tr8tJToJ0lMRrX
fpw5gp0mx05RIIVk80H66MpDnYHP8PkDOciGW89TukoKmm0i2sX6paY/BOFHYQ8F
+u5b+948HVfFmrhHTWaTgV34T3pdVt4lLhfZWcjZsdssEmg3wQQMAgH+39F5q2xp
3pVGDGHHvdA69D5dD4MuOzk40MD3QyTTH+2WbloFx9I5wBHKllvlfmGKlg1IGs2H
60nQPj5UG/WObBqbTzs6Nlu6RPubLQCVUeovu+DBLqn6jW21z7MybYESM/BD/ElF
/0GmBNTNkgdd81oWdJtjdf1gOKQjDEEWaReuPngDXf/h9eqGpUrJPo0eY2YBOG9+
hQtyq+raleBzXrEfBBYNC9FSrvp1TOtWTsrsyOkIansBlGzzuOWgZUY2jnHMUwyM
tqg6jDN620ixQtFeja0kFyeYKy89j8cvZle/GQik8+2vmOfu13VZDIe4uLDhS4ds
c9bSdiV5OSujWgiVpG0jEUEIZ/NyRpVSZpCYOYpDh1k3GZRqbinEBDC+Uun5X3u6
cTluoYo+KKi1uaiTI/hyNw1N9ZkhK7E9wjSSGT0Lhe9pacOXZdrf/PIzuxV68Cvd
fharvPK9jpsnzgdNH0VMJ+KMWDUxe4a490YBuXhdX+y8ZIa3akSc8KcBl/pgbE9p
xFrNaRrv/gNxDP82WvshhuqA5VSkftyTTpIm+UORcVC6WnanDHKzRM5BTRNWRqaQ
9j/Ax9GKA4bejojTR7PtUWULgVQcla0QEc+q7UAT4vhVUzY53YOKDn45rd6S8Xau
MbA1v0E0MBGo14gtPW9QN3g0XlfZkl1N+PGG8t7Fq4U6ZEuFj2GWJuzf7BbECxpB
LCSrZVLvZw6aHXR0itLtorHTXd7WIIWGBkGYc0qtqdZ+pwQIMZhfmO4W5V3O1xHm
vhm8+Usdh089GNY9h9KtsNMq98MeRwz/0jdAQa1dgRDE6RLvy0kWjF0m2+igYlZ8
261Pr+B2vZhoVdtA6ZDzuejWiiKQDuqpobU+JTmabfPdtOwzjxjU+/rrxR0yo8rz
Bt1ZGpIyuyeOUEnZJgNq5mcLy915Chbq97jSrZY3OqGbvaaSjaDpxLkf9S7SN7vi
r88XbP2CdoSc5Lbl0VCrDMGbFVCPrrtNYD04VBWkKDvOdecttbRSkSo9+x0cH+71
qUJKxGnz2EY04s/bcdNslCw80ac00JIl2LpPQHDCi/JRPdTFRpxLeiusByyqf9gG
rYKKzHZT6rpMnfFxNVFlRjgAe4L6YkcBAd1fqnqu94m82dTjcc5gY4py2Gmhw8Nx
rtw6Dg2vNEWX6ylHdbSBshbfQXeK9bFyacGXDZX/l7OV9zSt3OpZ0JvgLE+ac5lS
Td2GVjnKOHmzzMrAVKSYn5nXYYqg1Z1iW8vmBPh3tMf3VzkNaH0DO1ofaUD10Nok
cI/vflyziN3Q6NEk2uSNYGIYe7H9EBvuyAEQwfVnS5EwMoDlcUfL5K0XkJ2o8yF2
fyWI5a5A5BSQDM5mTSxV+bcH2jG7j37oMEwthKyz1KdywGMtlVlG3+NYJ+n+OM5K
GY24w0jJhRk97uzRTwEgRVpGj2+ENButqL7hsfIzDtm45Gltd/gxkjexpfTj6FXZ
pjL9/0Oczv+GuUkNOH0dt6kvQG7fbd1P85zbJ80+BqhU98VsyJKwHup78hQEQu2l
AREtnDjJxGVsWzvmE1x5oxB8FbYx3XkeXshvVLRvQKiBpqgvDNkFNh5/+dvcQbUw
N70aysEVGTdRxDDET4HXbRtQKOaTJVRTsrEP7gRSiwLEDyeYPGjJ0afVgJf7d6hd
0M0hncdb/XwSVqiSs8yz7FMRWmVAuxX8FJ7F97+ke6U/MRRKMcwncpzwfyNtBqSJ
pW3rDzCcb7PlZg23OFrfTmZH8MwHq0wErdmVZVqkWH1Bn0aLMqWbR6G7ob7ddSH+
rUbgtxqSjZ7xGvkNRJPjDtdyEcjqrKrQrh5PJwsRwjyPN6NC+NtxWlyuIoYZwL1+
15HV+bV1YjtEcSjV0CIzziISJwq81oS/jlAaG0z7+mOXfPKd0Jkg3L6BLZvudmbf
zBOQe3qA3xo6u58IhucTZvvkkxDyGAqsBDkrEe7+DZypT9wrNMw3NjWHQn5KmMJy
lUXDtgbk7BZMo0jC4kFcxo5KfJM1jmFDBEfF9RLp5WGOMMmAV+XEXOjiDQVUvKQ3
c6qh6dz15nbl4LBoYvMxTosfTgBEqWOqz0JONXLXH7ikMx/G1KgQG/Mf89YYHgSH
egj+uF8XQ+dzDsQLPvwC2jW6e672ThDSzT/N0phQk66Yeg2uKJ6GUalTmsCEAfyt
nJEDVnKXDMDOq7Rn/i/bZ5H4jvpdLqOP3w5VwVjUctFHQw1k0OAvbWqI+pT8XLgk
cZpm9MQbMIhnjh1OpkeuyKa4Rp6P8GN5JQJiQMHIlTQKRs5UhBlZyLdEcfcoWPN/
SeAP7aNU6yqfKdevdJE9w8u5KcsDsDY/WXxsySqRJAXH8jZrmW3qE+Jh/KT2/9lL
NRSfA4uutpL3Y3R5tEURk81xTDIjv54YuP9A6ymmF1tQVH5lpBJiKmE6VOWixbc7
o2QTDjI3pBO0BPRif8fFF77pVq3g/WQIly5zqR3Ff4JOXqd8nmeXU/OaAC5gsW2c
EEZ0Ak5+2vy9fIXXG3cwh92oCm5TpOQ3fBh7VrfioZv86qauNMavF5UpP3j3lL9O
lRSb5d/MwOsefq+OQD0+fwhK24a/+SuNwUhzoaTiYm8z6u2NIfFXF9aRCuATVdM+
0qL0HYxumP7yjYLo5grY/TCr/tnkDVqVsOR11x+mqsLApNKFNEr7ShN281TWuG4t
iN8Ioa/9oQWCjwZFM0Dj/VayMLgUXmANagUNIe7Jy2M6//QED+jRu+zFi4CT550F
RPpGNJo+eR0sp6/vREaLjdXz6Q1rYNnbv5BczvJHFNt9R508BbEGsAKrDvBFQWqN
hfsqrygJvSdhuzD0THV9FZqKqpoVXyfj81/6MINmoVdMoZCdqayffUp6VXMSz4cX
YYiAgbvbSmnecLfsrAfNSPCaIMtnQbttDdrOv1LWoJexx7VM6/tDO8NUhSnPA1/R
aFOF5ksmJuKdKMU1a7UeU6Hxq/NJvFUXmmY5Fj+LATJuNHYWw9xYlj8i+SFILb+k
Qr+tCSNRDf7e4goMv9xeh+axEHv3j3j2lpRRcQ/mSc5ewHCuQQJreSHfc/nMYSBi
NPjkanoVmDIkKUc4Z64Q6PrB3d0WDD8y8vwXvjhJtrX0LoSwDtrZnN6gza7Z72Cp
gpJ0gPHKIYFEO4Vugqc2i5l3WMLJB7Lnm/b9wX0sMSVqA7lLn5WFxhwh6Jv06Jku
dM7XuYm4uvvRewByWCuiMO8bWv9GT4AjfJL//NyeEYrU1I+n25dcXfCnZNqWdE2H
noZce1nqSTE/1LddN9bFKeKnHC3Z0kQ9DSRIiJgvvWMR3idjfnd0Rso4krnmxcjK
3aCl3R1gISqRS+2DjxcvQ0xt7OZbrkwCiasuqNzZajTVoqOfRX3OIrrx5XBcEJZf
HdbLvHfYYUc+wHwh6mA27yyfRpDOeAoKTuodkFx58J8fJTsUu+sMWKXcdY4p1/54
d2u/JAhQBjtMvC0YYFD5fqsnK4itVA+34oytRF0gUqbx4CYXQ51O2MPlEieTgyjz
opVlpIVx9GeiDcqFzbcsOn+z4NVuVTYwUvuL0286LkMNzE+6kLJ+8CRFvVkWsSXR
9N4Ms0E98aAFnAjYbGMClsHjQ5aNYF0Aq/U0I6M3IniRNac+r6rIVuxvZXW9B+yV
47nQnC/UvqjJp0ZtCzuKRpYL1Rg+DIrGoLfSroPw1j5GBLFF1OGk5uq5h1jBZtDu
2jc/FN1bPH5uXw+1e7HP2CcSlqAz4vb1oBu4FuYnHuSXGSFB2hd2qWQPOfya0/Z4
5dwc3yhVBn7WWEDWB7sIMLF3PjvnfyvmRGhhrX2TUU0hb8ZsFK11s4R8/76zySiw
gaJqpykSsTkUqEAsoJZMrEGKdYsjgnCca4Xt9DTALeq4jzLQ2Ncap71M27jQrpZl
LBj/8K7EkKMA17icmluXqmnCyLtkdHCxSrNp0xK/G+Zd9GLyprkWuZo065YsOBVL
rzF5Z2Zj8l5Iqo2Q2yMUMOhYNfMjWOpBgWRCkjdiI0HilCoAzFVZ8mwz41KBuRBL
k+y17Oytpfp+vAzQitm+rdSpiSfHtd4gcZrPN9OPOmW2GMRqap4tOhr9i+RTNOUW
zwnz79mYWxm+eB5NpWvq3I8JeUw0yK4Y38wnPiTkjZunO0cTNpJqBB2B4ajrL2Yf
4gFjmsO3py7RSvjKgUENewPcQuDe23zaO2EwR3gTaGXyL7MnWl7irepMOWuJWzrk
ewjkTG0iwfIbK9ULgAFvDnypIVXog9lc1HWBLIA5dRj148+WhCukCrXYV4GdY3sj
YfoQDihrfmmSYG6aqADDrlnJLTE2r8wG6vahvGCSoLG2NHWy3AvFwSvyrYPNu6vC
ukEGO2/CRug+PXrZLk2K9JoRnoB3jNxQxsMJmbfGHeTwUD2FK0HEU57XZmHzDmNU
jYVVEsGe239P2qgZpqCZfKauZUWZIXxKUz1mXr9XUJLGVOo83C0K4HciGNt5hh+9
LID1oB3oYWC0Yy3Ug33CeJISN7lZ9UXDji+SoBG6rz+wCrJ/Bnx67LQSmpQYduYU
hdTEDnJ9pcKwTCyBqxoNgRSdaQaSK7wtiB6XSlnNLQPoQIDi1Mp896yvshJgiNSO
0jOJXsAgLKDkaiUGG3AreFGTA2V2vaNoTcfxUMLzLgzzAFZzMDqDmFfjUfBOO8uo
FvK080EG86BIfEiYc1q3kmXxrw+cCyPEzmL0Hgf5QeWyVl8NXkEdMH1Q5KJo+hCU
F+lrRiT7lOiRU95Qm+pQmZ1AJG26jwNVdMydJhBuBuRXi5kHJejdAXFgvi539F0D
2gXRwL2OIm0xoo4tRjnyPV5cUD2DvNfEGfk8k7KVdd+hqwD5UhJtCRN5pZkDG2YC
ZglubtaSsO9p0si3qU1P0SNoSmwGRXEDE8R85iLoPYs7/u85d1scUz/FjRC7tM1f
6jqLuOZwkRjL9T9niCyNMJFWjxmXtK7jiSU+pM6d/i4GvitL6pt8G7xyyUvjX+gn
TvzisFty0sKfbkyCYBhfIiu7sWqPrVi28AjS0YwUD71L16RVAmr/KF3aI18N5nU1
JqlpBH9/CCkhetiD/8UP/yWetdCkutdi1NM0WOQtkN1Vjz7h/nrhY5CoRjZDJ7Sk
yFYZTdT9h1YOBSc5lg4hTCsFPfxm93qwGuPCwbEyMoHe0DEqlNeEDNSIAazZse94
BQDKY2Vgs6j5lqWfFo32g8M+ukv0rMYaOl/r2XE8TPdKU01ze/elK3ja+AEHVnAF
47h9idQYIqjsq7zdtTBLidF4muv3CfH/2nS+p+sc6SoYpL0RXJ2MBbNx/uExQmGe
iXuPR5RG5+apTxJ5BorZTGasiDBubDA6HSK0mcglLJEusdrt/cf2LxhjiUt+AL7s
7LD/vEq3zQ5NP09P3dN8V+TKP9XP292NzEeM9d6o6nMVU0476glrMo+liKcojjzD
KeQwmMDfaeP4Ppi0KTG29Nxt2xP+dFvH19keDM4iNskCTQ/ubTrhUxrvgwM/CY2S
3vKXYvnaIm6au4KF+GbwWtD2DaSi8KpF4QLoRKFOxzlC/5hi+KoZEIzNmEtfq/Jf
tUeK/JdgSb7ZuKw2CngqjgtGumzFwvtfJF+CA7T11q6zTqfABnyaO02blmMCLzpp
+Unkk8aOV2xhmb5WT2V8T1G8ZA9BpQaAzw3v7TDUlUQYuwEyBnSCZByxTrPtSaJQ
usE7FofbLmbhQNusVImX+FDTloIXp9gFEHE3wY2nY0Zr0iqdB2JMrzI6WiXynjmt
PbyLbdRFKzU5CevHhbfwgUohYeBI7buzUJRz7y3ty2eQPQjxCtJL4LGxCZYRhPCD
qkzgcOcpZWQqzu0Sie5JJ1cQ9t8H7Jen0fuz4s7nJO74iuvpaN/vWGxR4C7AycEC
vChHVuiN+eT/Eh8orESI7Q0vV5UCwm6fORepgr0KQgaZi+y8rxWAQfW5XHU8LolO
2QXeu0CraLhR9M0pPOnyH39IC2jqfycOx2lR6dtdFVeq6Vm3YeSUXDZvoOpnszDl
50EDSHiqu7vbETr+6muvtCTcsrqV0l6jo5m/729B7irYMlNOlaPqt9If0vAJKGD/
aKV1SM37P5rNSkFSOclr9JIX+vYOUepPoRgZHl9BREj5Aw+bEKXlpS7acZmOMkI0
GTd9ocHzktzeYF/8QDPnuJ4mMmZoXcGu3uWP5xqW4PKmuPHRGrBOvA5XyWOk3xXD
a1YmqV9uV3L6mqA/6u3ZwMkKGkyq7m2D4/o17U5AVEGvxMP7yZTxi3kFoPKM1NWS
Yj42+ehRv/PjijJU/m2MtVvy3yCSWRzi1gLPdPOCEf3qr4HuieTx4YU18kps63en
IKzvZL79Cft9r+bUjcDNuqb9KSqfKxjCE5YCdQYODP7LhKFnTIHKNFsqnj5UZ054
Ql4gnLG9o99/hLs/WRAsQQVdYKfpNKyA1N9xHfG5FQc9NdvX9F9TlQ6Rj9e2qyvV
WBdg8pnCv4tq44ZEBZp4ehjDPxQjT8m7jhHMz1CPsF2vNCWytoBZrqYikS9S4eSf
qu4vTiMOgTTl3nyOvEdwsmOoGcXzFAlNuBC6hcTEWOpdO7qxVT815FGv86hyr8qx
tcrHM1ZeXw//Go2gfHoe6jEgqchWZj34t/Hkgg4Cx+3I7IlXpsWgrkJyhrRwlgEQ
Stenu+dcQyljhifiw6FATnKVpzaU5TIpCmf2k7b6DKTb43QEBRcwLmAIHLqSkATb
8TTc0Eq+fOzeMG4Aqe5obxm0OvvfRIbWURSjQabgUgrZS4/HWvXxtkirksVsjRKC
IdFkPTprKlDccVa5f9Slu1i0+0+cv32Uex3kFb2/qAcurx677zAJ3vroSR0qGWN8
mUOfUFy5aA2BoIuCI4Ly3y346QuR+8go9KwlLTivyFMpOgw+n4poTl/1DtHLlYt3
sAdp+u/Y88wysOw2Q4vOvQUVKRKMLj4eQqlPjzcE8b5JqfrPPE5GIzq5sbK1KO/F
FxNEK4ii11QQe7gexdhtUQM/uDD5+DhjuvRmTtjlDi4Xz3WKAEEu5LxKPFFJNtn0
4ECtiXx/bnNINIAMIwx98eSVAUN5m9Lb8ugTG/Qc6h0B7M+RWu4b/vR9noy15pMJ
zxSaKvm2dgf8qoKlDVTPTcyR1H98v7/UeGS36n0n+e0VqU6PE+DVF+K+QKNDM05n
pbiquBTjp0Knki0lzdgZee7pvyYyKSb5TTCCNI+5SkVsDTN5ZpTrr6lzbKILvHtw
T31RyWAgvpa05j+qohlAYsRNsb+7f1Lz81PDuDtb0rrH0E/ofZ4WDyvvtRW0M9jD
zda09yf5SMCbTBW79W/9xloQ8Bqf4Ye4y/M/8YwVt8X/WnYAJBlFstd/kv0p2Xee
J79CjHI21goAsh3bv9TpYpVV8zQhN0a8xtUWqscYsh7T/9aF7sJyK4tK3Y+NdAfS
fBRzoGbFB7hMDxtiEwZ2QjliVT13OOlIh40I7Hy4kOUzlGd/A+nIq+lChZddOyZ4
NFlqPRr3zJJMCFHrgWzLhmb0WFR6esSClFqCb+mgLNYYubznN83h0oRX/FDICMzQ
NDiep72d/9g1G/3Q9iV/wxR+SWJGIrVnEjpBh7g8KkEmm2Rmh/idL/hzWZ+f1VDF
B4yBuyAezXMXnYp7v4pmn0jsI5ON+hJ26kBYtCCj11aY/vs8+eKbc4gn8XDMsbZv
8FO35VwXc2zoUQ67CZUfL3JVRMJUDVU7IX3Y+gexi80YNrAFi/d9yGHB1qiXZO3z
xi72JpkZiZaox/dUcPgj6ZyMhYRYGTvVxFNmmff6y1kBC+y2UR/+GkW8PmPOw/fj
Tgi8hqy+ekzh33qGlyQUvaGdZeGtnI5y4NV3pd8HAaZUx9TpZdJmjg47bEGd3ceB
o5gTVkUpSOTQAY0QTyr0Nnl6m41T4hYRfXCcCDkWwEEI4kkhbyYCMK9lTq75yeAT
cW/W2Yg2MPcJh4VHBFJ1b6Tj1fRxGr/sB9M0mEtBaSoY2pKAvwLaR5tUhwF+ivut
w60CdMpqLYvQ6RTucDNtE7Of0YCHqy0YFjwGrGuW2Rnjz4R1hCpEPgtuy0DQxNwH
rc/qHIAQrNVwlg8iXQtI8ijND+oOytn4/QRE8UbFIyFxJIFz40qMQt1vCwn258fC
chuRzVJNyMLzXJXZUODze3ktwjtGsx9m0U9gbFPAQpMZbfmhB6ssZygQ2d0yDlFW
1zXUe2MJG3JEGZykrP73vV4Nh5wRuwTw2vWajSHbMIcd2ARml+tSmYRLS6010741
oh6VAUHGbRhYZ4LCLZ1e8EzzPJfBHDgh056mCvt/NxAtn75I5ePhIXgT69L8YFoS
APDIxgHfGRdr9Guiu/dTmtlNWA+uOXdvgn6T52Dw0MKtKs7V3jQwKyu5Bvb+O98j
5Tt50Fa6a0wrT88d4waeU3YnL34GLXvrSF59NRcBNQQzktlDLzGJwc+n3+x34VZT
hX5U7YFkvGYk+wip9EYpmdkeuSOA/rYRwvPN1bJLdGvA472tG9YpBKYoeYSkZzwh
3AhV6EyR5r8reTGgrJDWbXWkme/NDcmFJ71CPoLEVwXLc9/5OYKzj/5J95dcQFDf
ZA8PQ+5hQRYOPYu02jK8VLl91tPbV7c44VxWNjErCGtOvBl/wm0ioIjmDAlVWx12
aKfX1jgSLjj/CPCCHE4I/v+s6hwseT25K6lvaAyMmzhBS0XKD5B3N0q5j/Ajj++0
Il/+MoR5BsR/c7LG+LfjZJ+j/M0DjSO3UOqkEUkaf5lrpWyAUozdshwYHrt1UMWT
fE0sliYXr3VDZIJ9Xgt8UDEn9AQUrDgjB9tZfFO9uypIOZOKteMYHJMSUzI142GZ
nMcR2pDxOQtVV2Rft5751I4dWSpM10hGtpLQScHsD56y22d9HpJ8MBchRtY22ron
W/aRpbBo8rsMXdkFngsPlBkQGVWzPNNI9+phAHI0tPeIfxRFqXx8cFE+aBbT0R3W
OmNnWBMQP8Uvi0C9JK/Hpq47XuCWXD4YzpuMo8LUGTDPZW3+Ers3wJETREeUvNKm
cRvgmAigtPgkjHsvdovM5rvzqiyASlGfotKBCs3yJRRmwWTbu9eFG9UODLgAuX3P
aOSXngALHlFbeMurIFqIjsuVk7xLDxCbYFdjsvL06aQ/E+ZY9G5F7mh8V8GhuID/
O+bAi2bRX2K/aP4jbnq+I3VTDB3MPbY262yYiVkenq05eIRpvt4hYRN/TcUo9lLA
ZY6XD3pPesjKtPbHqqVPjMkhb/9rC6hJCwzyp4feTkduZQyi07HIIrtAdjDW5JJ0
ciYdpKbNPQjwJs+tYld49SAp8nAqvlhrrh4QLcO0SOTWQ6WOul2xYvBgoHTh5n+V
jK6FkQQl/nIA+dbgSGOZLPvXatbazXcb6z4n8BmJgy2LSScWalpW24awu/boNbMU
RUEQAjPVs/JnFahCYRkZIaAJTaq3VvI6KSiYVtbXdT3EM0kE5fU3zUbWe5Cdeq/3
/LpxSxB1JcbM4xyDO6f9Oeam74s0T0jqpVdfRpi7qqwcKYA+V6dqO+Ch1O3907nT
uMH4dVAVu3yDNVO26bSD0El5XRedxP5upd/E7/vxC2NAiugG1paT3LddQT8QZXiA
bavNgUQxTZ0bDIhjSm+5Uigk+XDAWsfcQgplyY+9FtH4kTEuGmZWuSsOx4xCUL2h
AknxwRjS6yHLz1rEfruIuMioq8r4jey9wwgFmktISwcVFlCj3jf4a6CVa7SfLn29
L+R8YobRe4bIRKxUF7jDqGp3FrYWCrkaAdGlN/EGPSO1u4vjP5o/00EIS9/QMlWJ
UYiW9fYGhjB+DF//JJc9LaEr1T0Xeb+lE/D8ihATYUiQYEPCSeOUyOAqJgiN7hsN
xR33hihrYIlfj53YpFHd+GsG0be7KfeyZRs1xdIFynfNYe5UdR23dfQiiPlw1r50
tQHxO1rwnTOhl84o/qiwkvap8FhqrfNjNsR8frXiWRXMN8oqQsBMB4O/yNTgjs3H
lqlflaAmkOyzItyVU5rPoMYZeylu/XkSFuhJL+RA09yBGzBY+4W3BFnMtos2cVai
UJ1hLKGw/7HD8R0nObTL4UODMVEBgFBR3HSJHFguC8vgOrlUYymmZO8t75bEfKdh
oo5HNJYddcbC87mGWxqbHg8BwfpSo6IWFmamzrs1vryXsQEh4pSWdBFBpPawEwUu
EJm73AzUk57hlxLfrAE0uq6bfAYdvKByeinrd8LGQ8a2LNqGH/AGJ0ncQojYX3KI
p02oZ6V5Q2RvpXEyOi5zyZkpDa/QDVc6Ho0emobEvEvb+ZmpvrrFXf+wDs4Es4cF
p8ACDVMTb1vnIhZzee8T+tNubdT6Kyuk78sUv3jvkUPKuuQOVx7MwbopMOoe0aTc
xddViiEDfpvivOHlfgdY5L9RQ62c2H1nFwGjaRnhELT1KkNzelIcC3R8vY48ospX
RyX+dPLXZZ5vNxQ+BKnDkeLLG0z/3hDIT9iLJJJcKLc2JhdJzVJeKAEMQW7QwiF6
BQbNAyqUFFIqPMyjy3831pTV3LmtAZJWZIVpIpRtPWqN44G/7to5+Bh43Su6ztJS
KPLX0bx2AJedraOaESgdeFluhfTyj417RqVI3JCKo4XMjvehlbM/OtkgSf7/Bt6n
szxA6YRvd+WVHz05FHyuopSVStC/fuoQli4RPdsIPuF2+nztNwK/f7m6H1/iRvWp
cMHJIqRcYdT4717w525UsRbJdBi8xGhXH56pHfKzChAa5lhbM78JLSRh5Gdb/e3g
AIva1r7vgmja/HQVtmpAok8pa/rkVIHux7UOLp6N6SmsfpJM/+JzpF3SuWr99aVp
lrVslWjdS52yg/txUSNJAgWtjSCoMMIFG4/ZXxcV1nHM1II2DaExIwa7D8gh4iwt
N/aWhN5x/xKV4w2A26J5pNfir9f+t+AAQYf+PoZOD/Ls5GJ4YXHSaBSfCJyT2CYp
gzJU/KNgrFjFifk5jTJypAUixUfRwdREFsQObPN0/puAInJujAnp3/UZ5gx3kLDk
XOgG2Gk4tMT5dSgvtf8DdWTFixWJUk5Yg78F4eU+ofNCsunrk5NSK+yyUPHxf8TC
0PjONhB0IK1sDgnq5ClcDduIL6IfqEXcNngmK5HFaMKBhIDqBtkjuLgQcwjEXYK1
XQ7EsYhAiY6w7IZqY7a/xvXMNsAAFGo/KwaeQbS6PNdPwI7M9WuFn1KBrzh39FLf
PSMtgU4PtWrvG3r1WyLKrniGlUsYEeJee0z8dNjvuCM9Nb6lvSFqAN8mbVmZomGl
AYN0ZzM8GB/XuWJhaQhta7990nSkPxNAuGXOPcNs9zsY/+OVIUbkbHkqInE9XiQF
LF8KZZMuGTM+p1uyQ1sAJuTN85BrIkLN9RRdAaSdTmSVQ8x9xp/7JykjPBQh5e39
iPvVwszp6LTTilQ3VQnDzrryM9rzpFF0zQNJnklIjT9tssSJQvb6jTGVQ/JQC+nK
8R0r6FToQ7DL9nLvSH7G30Up3/xK1ELRXaLE0WLEE4Eig8jr1NcSSn2M1b8hzsOA
Rfgglb9YUV1qGQDfeWomChNCmhwhT/+GbX5C3oLuOk5L3K84cmolcsH6Bx1aO26I
F90ZMm+jCujlVbPm3zBl+vvt2Aj4/C8KTM8zVquMpU1wc9T6xybDyx/Lk5ZQFNv9
6jBGNqkwGk1X1NN7PYveHmuQ5iSzjobKX/RxYuh92ad5PIBM/9yoXTNsDQSOu4z2
240R4tAtet/suQ+kXtvJxhteCZjGFnkClVFtu3UBwHYLknBmAE1QACp8+TXYcbR2
a4qcfQvTEqTHoKPhlOK2KVEbvZ6wFwCvG8N+aTsWuTyU6htV5AjZMPvDL8dejLgk
+xaKGBd8mDZGcgbEsOe/YWEyYHd71Sce7Eae/qiTxTurxJp1zjeZtxsqFHv9mZfy
dcHE0Fw0UCf7q48Et8o98bsJgKAh1z6rqAGDijXPBs027mAbC/gtxY01tjPf6Vcw
I9n389MZVDj1sBYo6Szg2iVlj0+HxLdryphNfoYCvVbCm8lEsvWlZL+e9OALCSyo
uWr3hygbQ5mmBhbOJKWbI/8lk9QWsOV4CD+A/MDDpWh5t8R/V2AyCeO4ubuAhg2o
PsLpGf+fztY5fLIDuMdnO0Ky/Bahd5uZ9eaHASlWTyIqDrygT5IyzhOI3JwG3hp/
2Xpc5odWkLpwD+/dDEj2Mzxk4Jlb4TqGtrzDg6Gh36T3sBOFR7M/iRzNSmLfH1tA
/pV7SZxhhp5JxbptRZjfmJlCxhAhh27I9YIJNBkvIfA0xTT2GycLXPt65cpZqQYZ
M8/xBgz+RvcwpIdr8rONx3E/imGF6+utrjbHoNFBQo3MLwqqrq46uNXspWAqrbOA
e3wiklznd8Vwkwg1ntUhe548zcAwZzhBUZGwL3Z26PZodczcBrIiwAAz+gWIGX5g
6urQnPTzhM2r5UAr2HOdc89Sf6NbCuTSb3MDgHe3RZJgczgk03U7SKSYRmLODmaq
yKGktV/Cx/dVZi8l2qHkHl4bPiyWb9fHBaNDLrwC0aeort9kU7P4wfGKX4gZTRI+
BBtgYYzN/eeA2aauNJ2//+1I2OL8WaQRumJ3PVppwSMGxa3yqVUcpPUCOBJNE5zc
JJfSLuU3mMvynwKw3P4uBUj496RuWGkGtxu3t05DdI0gnRxin6upFVui1ob/llaN
+4qt5U7pMfSIbEAAApdGuVsIkXbQX0Eqnw14O5v5k7XVWwOwjnAYXdkUHIQ15NKf
gIIHS2RkpUj/6inouISohLexBpPy3vbVFEoq5UgClKi4dV1Q5sE/WauTxI4V7tHm
EQU1j/utSdkvHHcUAK10MI5DLVOdH1y1J6XJ0ekk9BYfMC8+52m4y8Sa1t0BF7pd
PJ4aNEariAzpTDm4kPLAHzYgwnkxqFX1xIuRRDDtaxnraenXmtJJQnTfULZY8ujE
ZmzNxsvPqssJoB2wwsySqS47Iw/QtNQbi/EaX63p7VYmz+fvDxuYg7kUBsmcVQsc
voHfq0sCJKZ9bH9PhfCSBeiuOvQ0UvMzJ6lWdgXDiKLcz5VoJfc7VJ79sHTdv6Dr
cmFilHyVLcKSw0Gb9rTmny2mGRYIAdOXMV0gjW83bmpAOyoJgdSPA2qOphc3l3FZ
Dp3XYp67D3R0qGTWFimd7DOJa3Iwq7UGYp1uEgF/xO0uN3eed4oTFXMnjq1+i0XD
64wFIQZZQUqJdRBxCQ8P2WPj8CDlxx41t9dsM1+nY++UJ5czR8w+8N/aXNR7Tqiz
EwQDiF+5bgrUghB5U0L+DDOVyQSw/pV/EEikb/c/wMqgQy2jG4IJq+S+2Q2dbkX/
lMDd82mRFZnLEL/eCGuXpVU/Lkb0kS5a8mV8L+URGrr21+I6hD4Iv8e/7bhVozwP
oi4vsv2xRJ4y0Y1rjicOVOfSkuetJWCLFAaJ9e1ldFG+o7k18W3zFHTk6n3hV3jQ
mCyYnlLtSyGwuXfK3iBfm1zWSkLYFrU6V4b8yojwtm8WBlULE9S3VAf0jKwEDuI2
j4cOG2B/KxoSdXz7lYJWmxVw+E6kUzbqNC2G+EfEEq9yjb+iQ6EF74C7yCZsYsOH
I5eGLx0hTS+k5V6yBrqK5NMINPvT2eH6Zc+4pTAy1J+xoFUXW4Uhp/imWsMiOdNC
op3HkUvuJ3Af5fHDTrz4IZpa5sXYQmEPiwhjL9y9BeHmIR1OfHVCXIwkUhMbaUV6
3V9/fYXVW9uKXbFDF490QrxTvGsTbD8sKOe3afJChkXgiBAEyJ4Wp9Z8WT+RjP/t
3uYybTckWJ3XNoHvphyJPTL16aaFFXil8k6wHtuABysSC/CGPGRvaEHN2jcs4RrV
2VAveefh1gKZmolf9oWeoQqVuIrzRJ0TC7C6ClXjWfQ1QpH86O57Whqxxew9zVJV
iZ/ewnW57uzkd+SGsvmg831skvqCMZA3j8Ide7W83Hs90f4mNcUq/5+Ltieuv5Oq
GShw8vXNXQF9VOyG8bd5l+BOstUZGeUuCX/O/kFqHfIBUXvh9qWkWz6SUL4xlStH
1Kh8gCJDvej+eyGKCuZqubedaRiQzhGjidKzHl0c7A8O9LgyReew/0G+IbrxPEzC
yko37XH8bRgjF/7dDpit4Cs47ZoYBNqAeTczFNPAXn4TZko16eiwHYYK9D5n9WtH
CNSKUWNklL2TIo7vvsqw3MbfXemeekb+oSY6sLJwiJGspIKIn+ywSELpntff6p6d
sRd5a61PI3Vs4fjcLAAUVQWzFN1ws3vlVz6/MUiBETPdwqZOUJaKScUHrLBaHwde
kbZUE7hzZdszZPBzKF5ud9CQDhsI2Lfxzltaxk/ZtDdQxQT6/RqHtxi30QYGD/dk
U6aYkh07zO/CfW0p4lB0iWrqAELn5eEvUwM35+IbCaNbRoVh4VcMDSi3+Hh22zLR
D8rSjWxCxzc8HoTrq2fl1g52oRK2j2I9AWtTEC95wHOU3ZM8HrPwERLaPU/BKKeK
kK0MrJH4GCPGSXpRTRthMe8nYWmaFdT9+PhnklHrIB9Gl6zlik5AK/7q9hw0reVB
pCqIkZZpLHGyGEfDxj/lZn5a7wkbrWMNgPNaegrjlAgF6u5ov4KsM/KguBDbLA6y
dn1aSdkjJqb45Atxq0RsZ6xXrkhFXtUTQdoAGhB6x8odZlvjX0ZKnwytUxOBMIms
DqZ5CdA9rdDZ8yQXTvyn4gcioIr8vMALgtU73RtxQk6rIhGi7Q0i3Sxvg4H+PZte
h5u0A5XPTZ4ipsfXmovfVHNsJwrj0tHH2vQgjl0DQYN/IqP99nNxNRy6P5cm4ZNI
RrgtXBj2Q6pI/LAYk5FkufmEajrvmtTzQ54lR+ug4GfcnMlTBaW+mouoMiZVjHKf
c8TMGeW+Jk+rdcX7W8ON32p/eVMb/h3QbqMgI8YhkvTESjiygVs/ALFfSjmzCFc/
1WZXg0EzktllqEo1fkjkgiB9ILgqYgqjUrDKfY6gnO+r4Hdre0mdnsT4IsU7MeGj
RoNB9lZM7J1Uh0IqO7yYnax2ldiTp+3WmWw3q+acpzP2Me5nopNCKk0XOvd7sMvF
m00b2mMyntcwH0bpMKJ8Lxdo+w8eOM4jLWy41NHFulg+gqjO+KsgAXLZRIU8xcqZ
ioV1DVmNpU6pietLktxW7xQfH4Rid9ejlKyLQxVP4X+ZrG3vCsGS0sHeuv1/5BFs
jmX9Y7oP3lu+4vD8eTJW/MEQHlIZ3CuNgxqczRrIC9/KSc/xY7IIdY/AO7++QW3q
YxxVX6TiZTWtv3k0knFidOFEEUisweC/EEaa2EZMVLRiB82AT9C66AhwVG2zcc5M
7M/JXTWWY6ex9W/Ia0XhwaxwlDD/HeRKhxfUn+zVBuhRg2PSJAcfGoapxrcRr43r
TaDZtES3uDOjjnyk0llMLZG0+R9Fbpsgorjs7y9axbgm2QebirmkdbVOiY+fqxGI
ofRThywY65uyclcbTyumntJLrPy7iKD1LfwFBKC12qQyIv14881j2IBAyMib9SEH
VAtHzFbvWkqDzVFns4lGGkluZzPgXC1UX4vsoQyeJeCGtVaUszhPSPC6tAf6nhp5
xq92fhjnt41JN6foGiJVHdM/7YAY4/rM+qBScC/4ZGkug09Fw2S03ZX+SZlm6J1A
4a0Thfz1Rz92cBAx7aIyaQ2vcXl6DO28dFM7a/+VgR6r3nunZpCg2UAqUiJkw4x9
/sUSWgot7MdQfjr+O+UkO6fRfTlXS49ONR3rw+RcQmzg3Yjc+AFzT5MwgIL4O4tN
yjgnK89xeINYa1Gd/vY8MdR8ZMAPMuHmhBnngLyS+JWsW0jkuDlzlP3o4HvjFV8a
jfTSDwddIWkzVg5DQ75bpioma1JzaZw6odMTLeY3v9vMXCKZGla5Lwk2PrCwgT13
BPM4+ypojLwdt4wGqjaS8wm5lFT8p2VCpj2iwHUwys078bGNWcByG7TRQITSxnft
sUUiwWzYzO7Z4yBIoGam4dfzC8pQtkmqBoN/FwfZ5Sbvs59vPTJJW4b9bhW1xG5J
AiXpQ2l1GciubcvRNA4Pi5RsfztGFvOjnL+dVwDvpCoMa8n6fPuIvqqxs9kiJtJX
WB+kqG8gRtK2fh7hjRSn2EYWB6HtzfRmQ8CSdf53kFjHuOMPjtD+nvXfpzPJV3SL
BznrjVBfGGtw0jXyzk6Hk0JrB4mtbOGBGpjotesT2EyEUzowMHoavPDTYRzYsG6X
e4iMD44afsa1djSKcVjpL/PNdWr4facJW7CT+DhcA94gJqnAg3GGC5hLzB+iPbeC
N8TrINbbCCseSFJ+Jxi49onh/VAlwfCqhIBKollPsh8lheeYeXPi+SMspmrQP711
LqVX3ueP5MKjG7Z06+3AOuLxT9cML9eCyfguQ71CQBBzgX9BXxK1X1ZNCjKC6hk4
TaiLidbsy5nUPMZ8vg88/+li3X2Bj3bRziCcT8nJGxjxfvXtGfwky7TXMEvJeBQz
NdZdPfei0BxFlPukNQTW1jhmnJheH1JOh35ABtSX1kTq2rlUsQaElO4ttJpD1qkU
pPRIxviHrjPvY5XTHbBdnRQ9JmMfStc8RUWMVb4raOD3gpGFSbQlkQatCcN4iEms
Kh9IwkPPkF8W9kUJnxQJsqk3LYVMVZ7LQTfClbqmGpDL7OH/oEvUhQUyJkAVXRtD
cBnBijqQbvYDn8G4r62MP7g5SxCA4GoiN8Xpl4ab702O6Stw4BBq6RdirDV+HVnS
Wp52HP9uVbLOlBJgcx1DKKu5aYenEK7n2sJcWpPTbQrFDMszmm48YrqrFKyTvFHO
AuKXH2JVOPCZl/U38AOevdx2lg5n2Windqn6ZRP7VSJTXxp4XRUTTUVVvB/swTWr
86+ot6gvdml9brIbloBpkJLdwQHfU6jFqVKGwGTL0oVK48BiaoKDTOiKvNtgTs/9
OnEcVaSh/GGh8oqGQHssLE6KVxa43WoA1nAooh2qIG4Gn391kv0hOuxkz1PgYnMS
eirXpMR4vjj2+NMhYg2EDRUAdQ2DkcL7LCKw0NzigEOR5pRpERruibfIYVFlkmm3
gvS6ByAUtggpnBBPO+YIT+hDxWO+v7+glWdR/5WRExGRD64Kx4QJ9QkKih9rY8wo
+7u3wWd+qHGvceHxtuujg590Di0GsoDq62EcbgArdE5huQBl4NUJge8SQYjnTURK
sFmr6UIf5X7QkY/FfrsNCkEbv8uJEKHp+nBfh1M1l1YqspBhxUsldDIPv+flVGk8
eHWUfeJ2J4Tgj1Pohvv1wBgFGlHWfdyyGyL0oP5ZCAJWOcIxPxhLzSToceaz043m
IsrQtaGuWgtPxsA/mKm2gfiZ5ah3Hm+DW9BRpDFcPxFh7Yl5qOAOQmmJg2TLL1yz
jc+zCP2bjXzYJ2kjqhUjNnGZNPUCEVRmdSVon5h1DAciDRAfV29eSsap4sHBq26j
u73h2kugrheXHQKFbHmoU2a96stvMvL0eOmm+AhMyCmuMVYovisJPb8m8wrxCHZf
pHTFAfzCNzZ2jxZbecctSfT+7+Tba+BMZr9DbMKRvvNmSerR7GmcyKGWvLvH9EwE
xmziEK+eTx8BI2MXbh24QV7xzuHbjDJ6lPieTzeRYwPSAi1hd43MoyzzIDTYs1Fr
c4m3W10WiJIetLLNpDJw8Aun1bH3q2saA3kmJ9LMRPHDy6WL3Fu1EHggxp1kj8kR
H87mYHx6dYL8CllmGp4oyC7kNdbysgaj8NYMYFCC5oJIIMND4dKoNZG5Z6I6SWCy
VdILrV/1ZK+zoZ6T4iBowtUBSprGijty6PW3YM5BtrF0LLcnMXc3VXh7VfuOM6q+
oQRkIR4qeuLOulIcRa8AWCwyP4LSVHuBr3FfohUEdavAoPFT8wAzy+55BmLmIrEv
iL72PBofg+WfU4mNb6+GyJkAFxJ4mhUv5bwdf4P7Lbna6yuUtWW1W+IydzCuZZq7
lwNvZVN0x8AsJR3GtTx2JcUkindcJbHYuW5gWOlu2BpRm/JRbJ6j8UkXqccCovjm
yAURQMuFdSqAsxBH2FCfXAyZ5Q9bdY5ptn7DLaNpamCP9VSanjeJVMK0eHCFOkGf
vVWc7JRhhb2tmltjpiy8KNr4qJ5wi62+wvDu8fYo5rQy6McDYkv7gjAefIxNcD6e
5bQ+7ucYXsqfEgEzQVxPP6P+CE0AnNcqIPSzW0Hubs6rJFZlSaLL5DF+fN3aXw0b
7oPmEIiOe6EoSpGcuWtvkbv10NvpHKYZPT2NnxbjkB34C2bf+obS6sjXoF1RO+NC
td+vbjRmYqPRxKaIfjR1ZFNM27abd4onXy35excLo0ZdbVeYA+3w48nf3u57fzJb
nkllbzMKmBpdzMO19TSh1OTaYv/Iry+TqmFovAhoN7dJNuWwf6AEKui2oc9tvfK9
meIlFD1clHUYKvo2wGDfUVU59zwKXABSsQKIF01s3VxRyhGd9qo/yTCQ7B/89nbF
F98Z+IudTDeVjfsIcR03XXtWgmi2b4xI0SQzc0sQP86uZAc/VXlUliZcYd5lBp1V
tZxAEmtjstMp9XySdq5fA6ZXe+5t4CVm0Mss3Q2rMMYL4yI4PRdI5wVqzT4wOszm
hLsm9uu/+hj3LWYC/I/6N3FFb5Fzb7zZUbk7mTTbFFV+Vx6WsHvwgtH14vaolKmU
Il78RwFEVu04sP1Ril+JXnyNixhtKeDxTrs+KmX+9CbOKF6P0VnzXRUiVvHoQ7rM
g/eQt/8OtZKiVZfYnKe+amskINNSRqgxAiD0BSqa7zVDB+ENe7RWBlKOeKFQi0eF
GHkcYe3dPZwc1EwpFKtn/PQE8F5I9dcUq1T/E42NYPdXxkPHff/mwQt2YjwQgzUC
l5fMphGgkMcdSeDlnfV2qG0gMKz+KaCRcCXTbRgA6m0wDdPi+A828BMxAv1RYuoO
nNlB2Q4264K6eZ2SWWAridoFd44O8JPQgBVq633yorKdHtjIFMXlH8CNRyGDkIv5
tma8V1GpIKGO13K6LXnq0jW5PYAcV/uXm8fHSGVlKYKJxyDZhZ2urkMslWlF9LZT
MUTcgkrq0beNHx6x/oXO8qT8NtdvKRokV5BOPA6bro1HNaaLVjwhFfppJs1Sk9Nn
ZZpfN3znJ8cjD/BzPQL3Mf1HJIkT0sTFFMiALbZndOF7kE7RVmEdMH58/dLiudBk
jFwINb2OuqXe07Ckgp0X0qFQzEJaA9OEsntd96jTgvQTjwmI1FFuQXr6TwsLLxy4
t+L5WboeXhVhTqtf+NRiPCr0EuT6hn3GPYLjqHJ2s4/EVVEzTOTNTe4Rg+mgC/AJ
amHOxVYKgjTpd64TT+cxJBtMz6lQNxkGbfzjMzHhFVQrUM14yFZREB5r6GPqrpcX
JNN6HVobP+54WndWpxisi46dv953XlbFjLHmmCmyrtVLtmewW4Vx4kuL2DCqf0s/
+Yr19KrnLDYEBMxM+lWpDsAoaFcyWYk7xxSva+ChLbUYzetnZdQenGm86nHa5USu
F+gAH3cEjbnWhsjkzo9nbCyK2V/BEpSlXSxA6B+8PJxOsMsxZawxhxI1Q5QzV08n
iM4ejxuyW44Y9nsoaiKp3FLpcjiB5jA+5VJ70/CuTNZvlsjpKx44Qfc8TzxpeS8v
VD09KxhQcKcRQmwjL6RcOQp4O3ziaROFDQuxtAeF0cPaCJB9pUvzQB9xjzV59RQQ
V8GHzFgZiQqeTNommLXb7Izz6LcbnLy9pnGuS6Xs8bFKexb5cvZi2LsrKXrlKWdu
Pp72WkbbE6g3ycgRg9YQ0sympVsardHA7sgP0Lg78n22+4xN/w4tIZX0Ulb8atQe
U465JOxXdbRaHwEDbbEh05Nrx1dEse0T5U49MY7Vbd6GwxUNmacf6+X+KMmKUJx4
poyXmwjz3Y880S0+t5elqY0FBiDKng/oltTPMm/ihsTfzQQM7qF08PfK5A4M8sxH
gRtphTO22PB4MQzH3ii9w8HwHl5+p+MPyya+7ousSo03uH/XwFvDkcjp/1RMXG9F
eD776oIvjJ5ul0GdetlC0Jl2vS0R/Mor21DVmEXeUd4JflNoF4viGfbuLpj/9yh5
JfPA+ZmhYIWeuXkHok1COZ+/Ae/JM3yC23Sb1yc9ekFEM4AkKFvfGfywZkg6ZoSu
HBP4UUiB2jf7nL/VMPcq/XA7qYBc1kC7YkZED5Fclf9/2yy/Ixyk+iTNi3pwqqBm
1L4CipoWM2L6hcgJDaYWuvVq69+2tcPwDaLDzo4AeKRWsy+iXpnWb6BUlfc6fZCM
CiDrJn+bnS+DHm4Jy6u3WkUK2PEgnJfh8hew5fCMD/wfWxBYpZpIZ+JcenwEHFQ+
1a3U0HBZbDnvH3ERNduz9609Yfx0P2TosnMMZjKEUnCtB5TVxyENQX5A8zgvpfPE
4r8qyznNJuMQg3WO3TCWnfc1i0CA18Upsjie8+YbUCkNnqSRSJWaDVQj1JcT7ds2
Zg6xw7ZtMUjnqpYyoiaAqSa9YoG8ZY9VdqirdZhBdD2a8CKUchDfOzRtGCNHM0ow
p5fKoAppvB4Ns8Ytt6u5Fel+DDSlCcybJx2dg+OVylqbYsg0PXnB8AvawPwROuUG
GYqw+VyhmMvvK99bFm/kyBQzPeLToJ5qj2umgK4q5jdtanyKYzZzRLHNKW4Os+/j
M0AGetlcYKukFJu12pPVQHZtqaYfZeBXnY/UCYEYbBF/6bnasQJ6Z//WQsjDR/+n
RoVDv24RjM4R/O51YKMjI5+cQeMrzQSGzWqdjZ+j9+/cEpAdVbur5/ZrZYubsHqJ
hVelu65rwgf6dTB67lKy7zfCD+x15sx+ck1ieYej7vWufFnJeCMHRao3RC1/GN1V
4JIb0d5LzCCTnyKnOAByybj05MdnK+Tow/XTd9G0lIaoyYnERoWS3LbQPyuoqe9l
e2GD4d5JvJfGK6MhwMvYao6T/+/l4VYha2p4wyiHNfrRVM9KBTGz0i2t2X1o+G2z
tWDhmjFes9BLCgwxqekukH8k2XgZDz7ETucePllrUUhRQE/Cw1O7k51Sz8BdGqg6
SBHXin/I6/ajIaDZMil3RIbjjgXpiUIKWyXF45ih6dq+FhbjnFrtNUUiHWApEz3l
rMeLtvUvYC77JCrJ0EAqlMwzb3+y1n/g0NtobEUbQR/Hd8SQsqyknwFzG+VuTnTT
Vmd1Q9xTZ8f82tMJxsjj8J27/h1/ChSUdsU9fKmAiBOTQaz1aS8OJr33AmloOG5j
aNz3oQYnxwzcADh89/6WQlFpSI5weBPDz7pmR99LsqhtUvlws61jfFl2S2UhkxC6
oQUFNLseJWJBcU4Ztg50rb8KbOSVE3IfOzub0ES3JUpdjrE4hKcawEO4bDu7oZS/
fJtNePaCcRtXN5bASyVI0C6zZAbSB0rPBOCEEsGIG4yfpogn9R2S5E28GEnhvr0Q
G2QIg4ErKFNC13eGzMlXORt37hwmy3Dn/ltl1HYEYVBx3dDFXAmAD3YaTs0eE7Vw
lnbevtQwh9cStn2zCdThf+wJ8Azv1PYoW/HKqnzr80bcs/o8kYkqX9NbHQnKdiCl
4gUpH4g4ICCO665lZrgfOrM5E0QJ4q+sU7uKMatEQd/7Mnqw/j5Z/rh6WEhSKvDk
qgC0eqMKrrRKDrNzwkDnYUMUtb80FL5XmkWq6mbi2sPvhH8VUtLm+OcAyCiMMYut
KTyBdb6RJBC1wUkjLkMpoqPUL9hrN5mzzsV+K/tcZ33HF1/Bjwr3dk60wP06z+gr
WPhF/JVuQFXqgCc4VvyYn8RSavemLqBK+U/Idqph2WIXNsJDv6smhq3C6zRH4tYL
FAd5ACCAFbkgR1/B4DGTiaS/Przus9C3xG7RaSCfLUFzHGa4BUKuqYy2vKELw15k
F/NLShFAUIAs0N4BClkXGDD3DmpYMas2kc2+3/soN9UGBgpWPfzn1u/J3kbNSlVZ
2Lt9a4+7JwDEX7kIhtN0Wgsa3paESaFYJan0V4tCYbTw1/rBcGHwY2grqqQbS6Qh
rGRoqUhEDxCVrz/+AzfpuDimxaSTWhSGL8wrKVP1d3wH5SPHN7xPSzPQOXbhzgXY
Eh/aaWJtiR/IpQkZXZC3cPH+kE4DETlMs2O7PgDdnA4abVMCtnFguvRUVEfjWQl7
A6+DBaFqvt5UKE0MKDQWAiJ8HxRUyZnZQojVzuoeAGMbSWihZZNX0UEbrfGiavmg
45HnJO4kanSYPtOIEdLkgJBsdWeJVVmcd6A1yA/N4acJVeuCc6GC/lYBEP0Pwr7r
qaNjh7TL6Ojnk6YnlmVXijXMhIB9xVFHHRC3wToQ36Ex6cM8pukraHDtDZ9Ki1QI
4Uhip4JIf2i+MqhJycmd7HmrdRn2zdB16sIoKuJ6rI8KL5spApao0uQBUvNv8FQJ
EC4WFVCfHRpIoIlT+hzegrmJZl120zEu/Gb5fQ5ZAt6D1zT1BzG8gZ3F+mWjnsMw
oIUe7WaE/yVw6Vq9vbfKtZVNTWdQ93wUr3v8LDQWgXQeF3NqT7cjyWhlF7F0c3Vx
rrmQSf5/tXZmUAdZ7Yn1Pa+S6qRX+QLwDW4re4MvjRZMjpUhU7iTY3ZRMZtV6fbf
pNL83yQvfuNGUsb6Sla/cFRCBT18gXbCI+0dX92j/MT75URm5NR0lDngPdDf7qX4
q6u2o3GljH6TF4pA5FBNOqYkcrbVY3hprrfg22QpjKHBqApTdAEHlsHbdXwmoUq4
Cd/lePxoWjz86/ye9W1Gj8YozSdvDH+7b/7OVaHaldQEOTRYtjsA2Fnp+H+k2NH9
gmYrTZsCTnOwvBmvSjBWvZ/Ugnqhi+AG5KhXcGx6iiFM5JWaQirBV0OYXVCdPjhL
A4O6RTPWzU+OW9j97JC2WZ/tJcnKzBtBqDxMLsZdw0GXl+E9O37mn+zGwFVG2jXx
XTK+DZj2zciVUCHStzLQ8PMYdDpUeaLfNOnve8Gzbm2w1jne3uxcoy0yQaPs87x9
SF4fSJIo1IpR/7KF52Z4U/uOBK9vr6Wxt/CdIIQAWvcteRFxu9MAT/roXVlc59Cr
dvPp43kGrMY1DCYgA444f5Xd0m4G4Ycyofy1pPgvAeW1dVIdpjoTRpeezaioWa4K
/hmNgza/Sjc9EwQdwP/JUsxQ6c0H0xt1GY9suvv+e5OLM/9qPvYNoRpkk3+5+fEe
a6biNG5TAZL/TU6fU2TW29t6tAahle9bMdVKnQix04K0PlrF0QGVzlR7721eoFHx
WIBt7MiEQqD6NlTS3+y4rnsJDX1DuFspb76CXmIJs5bB1xyGKhZbVjk4lIlYCh8y
EeH48D0Z9tNx20UX7Zfr0Ylt1GVsOYor2gPshtJ+SwOqXsn+yXct688c4EP00Nb8
t2U0TgTPh2yNED1Pn/3SYpMO1CbtHJHjKFhjrUJY8bndG8oZq5O5XFMo/rJOQREt
MKeHxFj4nRLpqFcHWsOxFJDmmi2GFWWe0hwDMVSNKz0VqbhFQ6HwFuOHt3pNzw2k
tK7hZzyg31zIBnq7kPlkKr3+ssKSGyZEBPretEVCZlpBFw6iJWvniEBXU+A7/p9W
l2VxB9QD6Y4psquG/ATkjwYI9IHkTp9F8MFet7mhS9W6n77ZhGiTuqtBA4FrGRrV
lOHfzvyq44gZpouY5kuU3gVTLrv71J36TUlv5GowYqNjKDtF+GoGJxALVg9HQpQN
qSym9ebPOSihI/bp0uVNk9EowE35pbS6otooBnmCf+5OU4ZYM0YFiUGgFXslc8Yp
0VTegPDkfLvqmfsl9Hh5gvxW+YKDWw3g7aa8D3oPKEUcaJ+4K6aB8Hd3d60OmUob
TNbJgASL+MdNm3bV8WJsixeXAXTLOJ0qvqi5vOa5bf5qn4p70JqMYTpW63WH6qvX
B8Tz7E1OsNqbvraGYJD7xavpsZYz0gqPWW9ig8eTZOLq1aoGkTbspdp8j5KXQW0N
jPRVgQARU5KKfr9VmzGRlpxjfl6GuQONKASOEO4OlVRd0DS13VKlYxXTyJ4Bi2M9
X+zjN6xMnNs5Nj8PRSUrwdeKrn+kEHaBQI9nJFlae0fsQ0gNAlrYTUga5Z8aaPTG
S6OQGvivb5TknNkLLEXRrv4dqAIIRrDJ0qnoRf85b5mYwHAbLCi1kr+xzoCBzO+w
rA0ZIVY/sUq8cpZ5OHTQK6ghcRw3oDEIMfSGZX0jYgeZUaftPebkkewP5KeLGDay
j22/jLUpKbmf7GXuhhUmecQCHnnHRPhQrNGNpUPDQ4QrAis+HXf4HciBE+W5rupG
pc5h9oDPh8UgTGUrp83fer0n1G+Zbj2bo+jLDiV3ZG9t0L0Xnc2keWRXmm/qOSW7
H2Fa7ZxemIP1DS4cDAmRpuUzluwXTPAvB6YwsV49QlJXIK9GN080QbuLYGxhvVku
phMJPLSon0gUOcpc14IB1e49q8GezYasjJM5rw0ZhBx2fkm6cGxqB54xE6tiVynB
U6sqfmDlNK1mXn81mgsnrlue6qMyXegQu4N88AG6TvjKFaEbyYIuCiL2QJML5cMX
jJxbZqX4BAWO09iL56hSGogHGKPCo7ugj3DHK05i2duvHfZ9XhB5N7bS728fJbYF
r8P/DJp/HR4a4qyB13rJPkx75XTQembO3bi40RfyROPUSLvcIspAYnF1+2GXkvX4
I1NcafDCaTRKfgXmtKLrSAINMH9w6Zc3t5UH4UbwfAu+lp4eYOhHpsXmetVDA37d
d4M3YEUJq5hVXab7O+UyjdqIW9Nj5u3QO+2oh+Sl0PSvIpya5oH9bE79egQ7lHwQ
ph2veDe0tPFTpGyoJQUM7ISHGpXT/g650PmXhterpuKxOMJXWcQCtdzuvUTHeeL3
Vd7xIiKcSmv13eGjs1/hsaEtiyhZzreMybZ8KjAdLkvcT0rE1zsPESROHANTkQla
jmyLeoNb3PDyBik6yZL/dO3o9C004PMh22ukIZOz+zj7QDrOPs8vemKEp23sa1et
DLg3zbNy17+LyhkCVx8uhqB2TQ19PhIw3nHfQaERYObTAzm0ml2x3fzTwCHnQeT2
eYfFFfIQ/AE5HakdRJTqOHkvcf72c3pn4MijyWCgukUvfJiLpkdGhsgg1JajikF2
US45JKm5DTftOc6pHpSjXrnBTdp66M8XzYiCdg9YnTqpF2mv1Zu/DsUGgl/Bmmmt
yRF6kx8xQ3ZXSbsznSRcyFueyxWbo9ACdTBfDqeb+HQXQTW6OR4N3FyIJlPUiA1A
uDw/GqqtQ8kPTCmY7RvA23uSZu6fRsE7qmbdB4pkPwspk3LSM6u5xALr+Sdu0OqS
c40Tz+8ho7CdMvf+kDzVDeUrL7YLlfsk4CWrxaHZd6SwZ7UKlS6x6zPN+5gih+Mo
SSZYXoiY1f22lj2rpxzOMfA3w/Lxv/gYPOYX8Ug14xmw0KfyfXe1WdRZO2CwjZW8
W7l2yfzhZuRRDCcD2MZ8/oR2h+yHPX5bseVRgAw5COEpFkQxBJNhFSGv1Bm2F9KZ
chkAKnfdunLk7AcrxBXJFIbwV3V3yXKF0edh/tZsg3TyczBFXHiWIBkfzgEsbQoU
RBQ26aMSvHD/f+Ryk+JFiAfOdm3c++TQAMSsfeR3j5goBTqNwn35yaeQjGQKg4w1
Xva8jYk8AywMJGC/FfEot8XMZlbcN2yBlChgET1/bDKbk0xRk+bpMLxBgaFPDqnU
0H9A+x4T5UCVHLwey855qGVjY/YbBhKUyqandkK/RaDW4z5f0FTwFmBZryTK4dMq
qQKNnTnvKFXp6Rr5SQ/ghfvcl1ZWwbODSTVeURTCWzBjhg7HaRBM6PrAU1mfFiPK
UCRYbvYxB8yGNoNzZIQm7Kf9c8zDZ8mDSwoYneBXRWtE/fgViCaS4z1guUeapXbC
8mgvGGQDz1x/6aNBiqMZD5FSXROTKSbOBVjdE0jeKCt6grlEWOHRo6WB8tKlqrOo
vzC7+jRT+mRsO49Ta826w0ebsxRVXP1xgMZTFURvhwNSmGIQDhzePMg1PVquC/5N
veSVOCe3jjPsnVx7JbVYcA0FmYaWJZ+d5+uMQKDFd/Ns3IK/ieMgt2Eg86TWelVP
bEgPSjiPM6fNeFlf50eosAIn+UqcBDyojbEcx5QOnfIlYsVerO8ftuqmKzmdnN3B
73gQjmnu+cWnxDh1FsRuhsHd1OyJaPmdFAAt2ujOltwHQx7bCNFt6xUhA6jpzVGi
7feDHXUF+Mkax1MWHNgKkTvEgA3J6TtwY8Re2nUQo6pxMycFK1VrFYqiyRPhe6HZ
UYHEcWavwchP5zyTRwDadAJ0d434ysLXpxbMAX46oY0=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TmKwJrETHhLzjAYQx9q68sOyVbiIWG9A3cR25890dV1rMybeAhjLXIvZIp0WiIqw
EDlgJsyS/4XjF+b9xPcaTaJXVwelB8/hTQWRv1DDRPBErdpsN2lFREKjndIutahR
RBP5qTQQYjWe7PLdQAZykNs3p5x/QGYpYKkEBFQOKES1q/p+JCF3L/Bc4/mxpiC0
H8mrECi5UABf1Vt1dRsNSah5cs4fxnGehKaSNGN8Bj+PF0nIpXfkUlO3Ky4Grz9m
GPaqMoOf46ySshdogmJLn/xHVsXr3g4y6+Izs+gvG6K8KfneIyzqEjsFkHQ72TZW
WY9ahHQdml3X+PN4Oq1qpw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2752 )
`pragma protect data_block
MifbSjyTTXl0f5NKBZlHbX/zC4v7TbuPoWHGrHNoJRDnRtkhfjZbmh5IV4SHiz7g
LSlnZIB3lpXHEnruOYu/zgQcRQu/Sdctx1jhasG2IUHm9Qp5Sz9u/l3oMTtV93rQ
waj1nARHAABrqUNCl6m+ybBjnOd4i1jr/SOp6R8TTIhxEMKf/B4d41+rv8F2Zn1a
sz9p6BczQvBbpeK74RKo0nsIsI0QQnf1anA2S+eAla6JPCb551/OGDi5xFTcmiGV
oa6YEqBxwLbfQ46htpvTuCRPtEiLgT93EwRN6db5hJaf44vd5q5dOI7cq1BkLsBM
D5TzfbZJr7n6Kgo4Ng74+WgKimRZSpus1lqKp34gT2BITTZgCvo6aOWWS1+BQMAz
uDjBJ6l4mEgk6GY7yT8TbcbeNoRCi87W//U3qHRs7NsbER1i7KOIhqRIn0q+RXxJ
R/rX7wntwAw32k9ReGt3pwgUzJDLRpitOMJkGcuppN7Ze/OpK6woXTifb+9k5tdB
noHbf58ZF/lkOLQC6ouThyzgbwQgUPLbD81wMx6EbcSqhJqbkgu521rhVggSB1P+
gzjqeHSv18wSl4GKXZVyt7R/AKqs6yexryVDXMYwQFueZfEb66NJuZra3fXJ5DbS
IXw6LwMyxCtgL4S3Yi2eCE6OgL5wU37KZLPCzRSxWD7+kom25yq1qyTg+bggweLT
Wzn8zhgOyWhUBLZZAHVgmxqGSBKerAB5mYJx+otSl68PWUJl36wAJg4EFYrQfh90
97cHR/0r8F+2pBWOLyS/gTbxcgc76PdrjjP4uKmS9Td4zv6EFD727K3nvvC2UYlh
KM6e81dLuH4dqz2/Y+HD5d3mjwh5IjbcDKN06pVlctbK6y9GLOUvxoLMpkHVkQoo
mSCsMc1wFJ6btYuwBuUpb/HNNv3Kwx1JvD+gaw8o3kd6FHvAgDsR89PjwTr0QvBO
sKU/e6fp0kdSp2MFnhdeuDmPQHu/qnaDU421HsdkSplxtnzispHE1Mmgi+ORzKhk
lTj6iuaGfiXuHTtpdNJCQVuvYbSexTQXjGXzpkJHuK1yq+kXz9ZAiRgd5cFISZLm
CB5WYzu2T0bCSXOc5voIjWHtugvg3HGLx17+h0n9F4LqiYJrPvPR8hQchxjKBxcO
+LMMfVkQqWa02wYn6zxjNGgS6AS+sLZ9pDkW3CFA6m+Bt3uSPJF3QUT49d0GoIfd
Ngjk+TKRsRpiOZ2ieDc6ALo4W6o54dKqXTqQgMrn6tUqYI9vylLuTB8HtoZ47Yh/
Iy/HxuYdXdOmickpvyjh+sKKNHWOuCTBL3VvFROcWuKYbIY/iH+YinTrUzMGNW14
SzxOhjI1Qw2nltOCLjZX6Io1c8pEDwhGvjBTMYT4NTd+Fy+4E6ZKqPZpZp+mfyyC
T4xHYQw1FGfrMuQk+Gh1hxJxW4zTPwDXz/ZOdTHgJ3RIZX+niMNd7pco66RxdV23
X+Kg5+aahT07hZbsNWSGt1zdBB5ic7czduS/cpfUEjoOM/nxoi0c3ohxn/SlUWod
w483yNpZJA8nx9xl5I1pvnjY3TNiXNU5QxQ2bOgaWcULeCrd9EZodgKcqplhJxOQ
1P6avoQ1NX7hV9/KOacv6TU0I7Q1P3rE9M2j1LVel43Nx2Pf+vBTiYlou+Tt4FJO
PcI5uOQ9dNQuy5z/L8xHikyLSuQ8n27jJQquOz41kFMaF7659VIsaaGE3EyHTiSi
nCZQKwjgqhnmR8ap5RxI/K0xMX6Szq2bLok/ujZtTca6ZgbF2IdKmsJlxlZBXQWP
T/6xky1Gz6DwoqpPgKvi7aLLEWF2Ple0SpX0hfCXpbwwX1gV90LtrGOcdmaU7C0v
m1ip5DD6a714kALypc4qh5ETR/wsc4bKF3WYOnK/XwOqu3KoFLtrmjhvI8RrkCca
3H8vsuKLZI9lqrOpgz2HfsZTRYLwcfWYM2I1KWJvZV2LVKmLxsODrR/6DNabzjPH
eaSv8RM29X/Hm9n7vH+b7gY8ItdmqC3bnblU4tAqrKPXmjOtdY5I20hHerR1n0w7
0Gt6GvHqT7IOf1LQGOMM5QNSHExjBssFrVIUymryrkr1gGjqcBf8S/MMimAd8tIp
+zSyxE03IbjBGzNTF2uXbCT1JiDifRAIS3/BrVkE1Smoh/lUebXwKXV5Y+JO3ieo
oBAxSudJEBoEUe+vfnLoh36CcHo7nMz9S4kxlDPQSqRbmkQzRV9Wm69cddlTRvcM
NXz4vkl7G+JKJiv+U8n7ZoK/5UZJrtZPvIGIhp3f+gg+PXYahQb8dl4hYQcWHAgw
EzP7NkrD7lLis7m7ryQftRn1zr1moWlovY79uBn1zwL8YI8Zlm7ZyOPASWMr5hEx
UPIGcnkzzeL9MHZr2eXM6HWheEl3vB2P19nVwxhG/GtKqiGulRUeQ+6xCukCCZlQ
gGDT8YiZBZHhUl1BaF2w78e9b24h9cWKq3D0Sv32nltUYrelb6b5FJ6SLNxHF3nh
sLU1nJ94TBNEB6N3Ja9vdF4tMEy6RLy/HRWxXwqx0q1q6TtV+sVbkiYrGfXxNFj/
wYuxjgmAT5eyQ1KWKKEjp35QhukV0wAK+WFGbapZ+QfYwkYSqFYCRhKcjlFGNfWA
FRLBLbxT8tBPtnU/69dFdqYPGvA5ofJPB0X8HP/yQP9x0xKmi24+ILkiA+adH6NJ
Km9WBB4Jplo220PQlEv7ny7aZTAzBZGUTn50g/iFOtmkmFnsCTMOKpvqB/UM4dfM
Kn5oee4CSQJEV5EB7Fsk6zj+gfQQoFlA94OHBxRkN0t916J2/RCgTd/NPqKzFIwT
0LLGGrUOkVUTPNqEe2c1XXW4jMofusRFKDFfBDkDyYxAC+aOp+TMOmDHvA6ET3R3
EFc+gSfQPnv4R6PYhPyiTpfUf2R9ARSfOdgJK7c0FHO22O3tkJJIK4dnG/bq0KlD
hm4V2yTAPsPlZGyPM+VZhWPKRY7Jy6XU4l5LR3DmR8pTSZxekDeKGZP4XVug9y0n
zKrFPI72b7uI/tDS7MfobnEOnbpH5mx2JnD8H9BhAJ7Aa0NeZA5guLWPbXH/6r2k
pbWTl7bX1blBhvBjSzVyrGcxtXLEJp2tmWKxtrIKQg590NSCa0RZUla1Vwi7amsi
5L9reybHFL6s9xEmOU63GxikzEaakKrBBPJmUisyx7xCLbiF/Cq8hHNiCK3zKnpX
nJIfNvcoKCXBllr+MbJwciu7A5vvxWPycX0BboBAGYalcehfNrLHieg/2EbBM4Gx
1jVkr14haGAltvD5iNCnKJN0qx7hSkbU7OFctulkeWFcXlMKVgbjDUsc3i2fWwTQ
lTRvMcRo04rZpuMbp0swqrNgxI2nQbRIkzU0KkKwA3OKug59TNeft/PRub97Ecii
I6xeeLLuMg4xmqXvNjgDX3zjoZRBsJRCZOoDkIcK96DuKVZkXi3xHN8tZwohJFwB
CgDvmAZmhAjmEH9zAU2DKYw581DUTsXGiyGX37HIQVPJpC7VK4HVkRxcKpeLGB7u
jLkpzTpulIEmZc55HBt+FWg9wYPK1YvvjKyYnWU5lcp/YbyKrPWEfU94DTCZ8Evv
OHzOaFoc+AzQdZO+X9mIU2vydZLPRgk5Ac1C3LYq6rACFbgheo/XHlBY1d/D3PmN
fx1409geOaZ4DBuxO9rCVg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
QmgB2GqqB++C1ZD30QcCh5xXmVNRDxpzHwffOmlo9uuEErIRVIz67Ap2i2KvyS/1
h3Tj7OTconl7tUj/3iGztSQT7AJqeHsqR9Sbe/hLJ0k84z1SCbptltTPd6z0U2eP
M6NfRJkheCHwHOLxfB2sn0tteuHJaWIiY5QAhNtz/I2McPLVN7CRzjynPhTV4fKP
/ZNrJevOUXy5jIAlWF8y5atbVLO+Okw5vNKGeVfkejq5bchUC+rMQrw6te6ocWIN
9pov5NcRKVkZnYuy5UTy9cRRh7nW6xEO6NUmeXJOJmaEgyPfqLukmIBDLQaizflp
iKTGkr3SG1STcUJ31dRVUw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1824 )
`pragma protect data_block
fv/Ay1iDJ76SqooOjXO8OPzaTQs6zJfcIXm3VM+GsKIMW9Wzhk63nFQJLUMb9G1F
OJw2XqTg9hlwcji1oGMe4+5dnO6+j9bZlJcQ9RhKBeDtovyUMXkLv01IH7i00kyr
wuyVSKBggVsDzNqkgHKdU+I+pokckyLJufEvpmmqdBU75i3YPRjTVXHrk9czS9e2
PbOH3Hqho4DxyelIJR3yiZSlSGCXfXLZNNB+QGU8uKJ1avPN1F2uAk90TjEYAAel
rOALHiZDKj3/M2uxBHYdrbD/8sIhKxpBRVfQZd6rVTy+ayudOBO8jA9xyTkgOrjC
3ZrEYZBCNbzOzeONVwPtci0JB7vw15tvkooUKyItiFxQpbucW1dolx3j9mOjJwNh
/qf3y2bF0H7SjKhac4TM1TYVgK45Hy3JUHGnDMsxBieE6Hcre13cVTgTJLhLNsKF
3C5XasIWWHmK03L0nDh47F7G8Mivo9zEhPUib+TdUAGiojjbzpyBBNSrZv3F6HCY
cMhPeP/7JQZnARYj03SI3ddkFV0a9jMPHBrHUBykbFif/qr5mCklJ2X/e+DFgzcY
grKQO5+vCYoerb9gUM/SodsEyLSVor3AMZ7ZAZTOD85jBDuQvoO3/yf9jhhvLwRj
sSns3V8WOh3bRXv2YrhGOhMCv/3d0E8GEMJESoLSAAIbTg64BUuSEkihKYgUlMDl
F/RmGHQep8kYSAvGJS0bvdELaQ/QQtUny5idPWy9fgBrZuR73Kiwg1wJreDhG4x4
wcjtw3q3+t9SKE1VPdLydbtfiI2gGFQk2TgCmnoQjbXMZKlZKbfac6Ef5Z5UxSQh
HmEm86y7S8XzEq5YPu8aEWjF8rX6FsuQVduQwR6JoMp0QwqT4UUljMye/VOLjzhs
RinhHh7EXRLA0679y/DoXJN7rKnQdxahP6ZPPVu+ACHKp++wylLVHIlSfvQsl7PT
Rb/LaNDRHtyZ4/CN+EviEGtAlAALdf0DVhbAI50YN46fkeACZT/SLc8rN65d/JF4
/k5IZg18Px8zTnCImG6gIGqEYdQucJUhJnMYtLdMDaV9/aV1uSPiyuZ1UvKHWvFn
Id/e6X9fXE+R7xKLjJ8czBs03Z7iQfcQ4KY6D0jjOjxjCwZTNEuOyZDOiJITINP/
lqeVR7APd5o61ze9iwBGO3NsOzItjSaI8pGhkZ+bd3weSZe9aXYrPE/opaME9lBo
VvX6uvBP1auF19rhuclC7IcH4XBt4+bMxbk67HS9JFFFddzFrQCYAtewoARzHK1g
vS6gDezGDo1wwO9GUZkr1dombLo4VBd+GSRw5ooRtGdzfXcqUeT8H0xZ4ooS2xoG
FGuDkdpjSqMLW8bi1F23/C8rsHdpQu6GqBLs8AnCWqZebi/R40nVwCJa3TVKNd1S
PYMSB4dollDg4Oqlskq25faJZ0icR18o3MLbvxcEZTyWNhw+n9pYUV+B+ZnAnTff
pxNc61a6MMlIuGPSnSOOrTRwJne+SwrMeuMvofS8o5WWhvxLcA08+0Qcq1XnyPwy
i4MnArhmlN3LnT3410fS8WRpVafYzXrBO5gxeTiVmN5Xuga7AUNIMtMeishQ6CT7
gpCzq6/Sy2uTDxQ4lHs5t+BWr4kEJ7/tFhEwBN4G4MhPDaxBhatTYpbHDh1C8T06
xRMbhTu0VTy2ffMAiuMcU63dgv/tUHQ8hofRtKUXnIXxD2CoPJuoGv9/J7FkR5pd
ns+slRjgW3ieI0BbNSQGJxxn86RnVnloMcGX3xlLOJFkOHnOcL8K65lMwryv351x
Yvv9fU6rBB83pZwLBdx+p3MQoZxJZ0Iptl/gNVldtavNi054t2GwlKUOT3KO2SNh
R1oS8V9Tqr0SbPq4woqt8Ja3rIE/MyC+Vq+UjTIhGKtaDtZDk+Y761wfy3NdDr7K
dpOoljIM+dgr3WNwzdDgFFVyImNOLzSaCvB+pl+Eny4gbme0W2l8Bs/P26xw9geJ
B+8l3V9KY5Sve9ZO3lIj7obKMDNbBYt9txD9ewP83PkkQ/EEGoxSbDB9+1pN8qY/
KG9HQOej5eYiOyySMfw/yvxcljffNeIBdSPKPPi3f/Hk1CNJDerjI+S8ig2MS/qr
8pLnbOWcczI+wJaaaeV9416pjDziQqzy/d3qgMp33bgQNnpNjbr7YhPzhUxRziYp
6e5N9dPCG8Uut6dCU9ow3GM/LEfOxZO7zdkdPCCp+Jy0rV8NSEqHUCulIFQYskEz
2EwSmS1zgl0EeUxDNIDrTJPf5p7Gz7/kXoVT1zmvh5WamipxSua1SPrGRVYrcOAd
LYGnUuNch1jKMHE7xcXjKtKGeQp+J8II5ACqkat33/V/8jLfDp4dhCpH+TD7rvsF
6zAxJP2FWIdemedVsshfC4vTygo+hSxOpUS22L7B9MNOidK8KZSQARMXvA05/Cd9
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
U4p/+q3NoY8LmYmsTx/7226RT4NUx1yZEir/DjEMOSuVCB1ydC9g5an6NEbLxtEZ
LPzkmaGfDRiOkcXgJpksZyMdj/pAzbzHsWu0oWw19xX5wXhHn4/xXB54TKJ/ndrJ
6glG7nfsJKT78X6vRn0ZZBFKJJwGnrtLa4gfgPNL4Fr/XyHSIEEZmlg8DigRyo6d
cqtxuzBkxDAe2/XDoObXqmWMSyer71xWl2+75eiSH3yBMj4RR+HAyKJxyWm/N3a7
zGQCo4rCtHORmrRxhs/COQJ4xWcBNN6q76mKFlzjA5B8rxSRvgyENFRBo1TSf08X
fc6KiLAvkeWRKU1V7pEFHA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 57568 )
`pragma protect data_block
Yq5dm3oGBWPy0b9FI2YrUlr7Q4bN7inyycSeG/ReNntXSHvqd1UqV+JrtYa4di5n
OxF5gibFYTGPkV2QKJVWkV/gyBETaxeivjwowEcJ50tiCopkrwjMg/NyyquhnbRu
3sOTwCOtwAjuQsnReEfHkeCIUXffuB1sztgqUoXthAwwBnTvhP4G0y9IyN2m+ggZ
/H2Wz76EojsN2jbxFjULAnNsFgNTs1ZS5h2CJeNbTB7/b6hPwKm3w72wzr3VCubR
vIEg7NDuuR0MuN6JqmqiB5W+iVpLzHHaSe6nEPLrZCN7zoDa72BqIoc/4OAhSLpa
EuOfJTwei2pq3yYvlgM/Z4jO8bSnCUStsLl2kLZ4SKJvu9qdvwNYcNolJYTdNDM9
qR3IF17xuCN50J53XfFLFzv4AtL/VPgGBbr35Xw/RskEIYCaQZPcxVeQtMSXuM3k
2Em6dCXW6mD1j8+3xxjDy4lfOC4plnB9zDSmlCcVPB47cs1c/1HemXHsKSP4VVvO
SApWKTlw7zmPyU+iC3PiwUCvUxvcZhSKO05KH4waMwnuTJcPMwpZM7hWClDj4ZhI
U2Q8YtvG+9BdPMhPfpUcYi4CwuAilry0wXyIgX1/+NVsISvMJ6NHOEimWo+Aye+l
SNBpHROY2JyuJcBEbabGHrPyFesANe+B1I6YcdJ4zjzUNa1lX1HJe6L6IVUkw7/H
NnIG95qlW71sBox4+2hhl8qHXp2F2IOOBYpzxF57FlGz3Jq+Q6UTClrnC+DR0F+r
jmB+3iaxfAIeOrHMtnjybQrVII0getmBWpjB/GlkljB/NpRGpTzqFXDnSLIwDYiS
zSJaHhxe4sts1rMgGCNPym4mK5ilVeobKq/0X11bwXuSzLrizf4voKTxNjp8QN4K
JTb8VtoEVfXAF8f+Z/+HELip7CHNKXyI9Fm43drQTyQdtlhIFyzZurO7sDKix0gs
4DF14ek8vnqkUP/AZ/cs4yN3g5PuJ9dGPr3Y5J+Cw8h9x0d+M5XchnvVIm34OihN
ND84/WBVpqgWtw2Xfr56OZA3iBNzxOm/K0pnhEnvKPzX6wUkte+p3OhBmB9ps17i
nuSRDMcZLaSMgfQI0H0T6j00uttNq9RP6pYFAjGMh1uIZ3lZ79c/EWh6Aq7wpAJp
IYgbMAbSiFTniQPPTrcS9ab4t6m6CgqSGH0Qm+Pvbo9MLjFML4G0JYRJnfxaSFNo
a42zXOFarYybusfZ9KHEzvOS17ZQi+nF6kGIJTvQ4qvrWLakt3EdrvSLCxtvsQgX
Xnn4j7tdm70CuHaIX9h0n2JPpFVGuCxWy2F9LUZTfs9JMyUOEmxvufmEPJCQh/yb
GedA3hr72Oi8Y2zUK+PvK0zYDgd8osha3Yf5bkxMJqDi0cP0omeJH2Pmy+8rw8d2
ToL8gKFdYSN+ZAKoo/Q9vQmyQ3vV9/Qv49WpsNLNQUKFQ07qEg+joTn7DA/kFfki
HgCp9s8W5A+tahJFloqk5e/KIlE5fF5sEipSI99WvgkqZhWFKOBbLlDDbyjw/Fln
/elboXLAbX82DJBBZXlS3WJY80MaxfgvdvhXdZmPx6mA8M/Y8cch8gY1dQy3DtON
ntb9jhHyhoDLD7WK95q/SegwCLIdoEZ4RuoToRWTGEYMkykrtbRwt0o82ZO05d3n
nBxMeMydZx0nbxsMEnUFdAa4zN0v3kPjZi7hSrJXgrtpPwPwaXzpfuNZHAC1zVnN
H8ObNGF4OA3v4B22cbtu14FhDSBdeSuBek7+89LXQfEHc7sdKTz61V7ZY5Dw77fT
F3M55Uy7U8oz3rs57vCE4emm00qJspscxLaDT6+5nYStYLzILXR4izzrA+jA/yOI
pm5bx7NRLZi9c+JDjelHZUjjE0lEDYzEt4KglOhh1Zov8o6kWctvgxt+TVR+czNx
0GNDwoK867GdosjOq6u/+gPsoboDA/w7i/KDUEg3gCpyAYECO/LnrmqjXxPxg0NN
YoMbDXHjPt0GMLnC1zcnJrsUrsis+cmFkLuynEMEG4vA7UG5lCiVm0bnICxHQQir
dw1huSg04Bg5WzpZnd7DlIbZlDs1g6nHPwO+SH4UxV7HPvLFycCsxVN+eReRUnBO
KqJUgPzxiBWWhiEfem/8ezLXwDdG1B/Cf7rhfQfDN5B/DZrT8/RgCxq5AOXvVYr3
yEWraq7o1FJ8odhX1hpNPDBiEdmgZxXsnG8aDsZeP+w7wjFizsvrf09dysV0DgaP
KuNTbpjJXNu/H6y0UEw4//w55dIVvbCFrxd/RR6N2DjH0lsf3/p3lWFLWY5KzO6U
VW9pg89O9X4N4G2wNK63UGRoQbuxtJDKJWk/Gyv89GwB35HzhS4OS/uglef/Tf/X
eJNkrNcNRbl9MLfjp8ruQ1oc7elLSNzO+3Rjfpe9jRof4o6lcLS1UdDVa4FckGWm
sCARcfi/GsJo4lJCbemsbQ5eTcICE1+XLrxl+DWVxixPC1mJn72QE6k2QvAYJJlA
EqmenPiZ+dTxKM7rBLmpm/KlJyroPDS71kDvi94I6xTdDDU2iaRZKYa1gmCfybnu
WYW8GNPdSCoayd96Kd9zaRD1gyx/W8o339abLhtV1dkNLNoZ6cFbDNCAuIr/jBTP
pU7PBIa6DQwbGpaCLHtkcChA5q6AtElqBCa1pyFGWPdERGz1igp+t+znY1UAvxAT
n/Wys7MzDFLu17+HNSa0vgB3OUc8AnEZTxdfCzMq3TA+X2pU/aLXzuDu2j1qoVJt
bZje+jQmRmOfY5czI8mXBmFBk87WsQLaEFMa0BkJg7RwlYAf25ssw9/ECBfCgNjn
tQlUsIZ0LPFHFrBUPvLeUY5dRYG4r9A0qPYKIL048ec9ZUdbt/SGNC+pJYMGAZ48
0bL2Yj4BllyNhoWlpbvjIh5DMh+ordPaJz9OMUwl032z49y49DWaKikz2UeFkEEJ
QpuT9xmV9N1yG/DHhmzUgZz++N3JIwj5KAHJ55rBRajU2sHy7vTy8U8SVDFLSiYy
yIfcgkvOvFUWdtSW3TuHdzqg0ULJgiENxtPVaYgqkCM+3SMHx+YCaaInxzAQcmzA
phwnIXbcPe+IvaPCPmPmGqtBB1aYI+7F3WsQU4xDIRhH5XCTni8uncosozHdqi/D
du3tToydk5FDGlrF/PqkJqrAGnsZW5ZTP3GqSdo6SfOfq9OJRtEITsrXfoNI0qWg
HSMs3oAO8HJVi3vGT2uqohNAwYdN+sn1fuWaEl0Axqkgi+bel4VJCjkazJ+DZ1K6
/Hf1uRHKRYVGRulZpDFvk8c214s4HVNyIHQQGWGC7dl4g13GmPACgl4tC2Spzg5K
JIIpGWVPrYtOL/4NeTjLpwsscfP7qRFkAx+BtoKoRiK/7FkhR87xhWxg0ITxSf5R
z5jaq5DWLLfIbRR1riyMS+N44xcULwWsEzCSAbYg2ZgeEMdvnIx+Ae9pdvrQtYPj
ruazLWEgJQU07kIbMCazDH8sn5qnQD89fiBnSJixD1Nk8iGCDZT0i/+RpV7+LQPU
L4SuEaT1OomcTyEE9ah/Au6RJg1nEJpI8PsTkGjwcT3CuWk4xzb9SphFPjxXZslH
NmgK9bnT4ihX4bwf1udBwqPbXsUMrRlOOV2b4mwR4oITM9ZEPDgl/t6y8dKuWzOv
WXbSpNvkXWldzGvostpe3lj71VOFqXQjnzZx9WdnfqXbp7t0PTnXJ9BMUTTXnuK3
sLM7UpUG29rt7Bsaz2aUW/YjzxrUMGFN4FMIuZOQZUTaiSxDlidS0czQF6DjSWxx
VlTTbO+snXTbmT73+kozic1RWISaO4sOLgujjPk5Jz4uqeBM2Jwg0A2gI7k15FTR
w4uFTVKT1Xi/pKs7+4FORADN2KGpmUmJvQa4J0p6Ksc8CUVhrwIsxRA/BRx6W21k
qS0kyu3Nf8/gevTsCJBp4RPZg6Xq1WIrQTjMqZRJIuAP8DkR9413ZXWzo/13GKm5
KFP1HbXZrdUGnlEx3vQU85/XCIxPBPGyC+36kExGzTwN3Z5606pOfLKbO5YBuVxU
IfcGaz1v/3oGr0rDYgKzJvtANXHMvu8CVC3K/5nUd2zfGFSc9iDWJNrOa9HqBc/s
N9VM+UhfwWvslVYoMSTflkSE/xqBbDD8Q2zgDvEge+NZWgDJfcJ6sUAiGKwm9bTu
oApk4RcUfH071ScP3bZTDKmjs2H5VdpfXhaA0arlYesWySBLuGh5BylPES9bJNO9
Tj8HIlohTGiLbfYbuV1KM+Mc6eld0HEl1eqqrYSKAyusO7nIULP6cYWs90UqA/fs
UwN20+uZFMvYuXllZPTCmzzeczVJRO/7t99QwA9w3SQR8IH9A1s+5bQTyZpHTo7U
WSc4HuNfUC5cC92dtq3gUanhKnJTO3mwzK5MMM3waM932KJQEY/nrk4FlA4E3SeM
FySP3TBGqvXjXKLQHRBMvRGFkki9ERLy7GKtN2/ehqvMNeRVCmrKXQOb2SaTpOOP
8+PbPy70DNdFZhEnt9StWMmXUva5+mbZcndrDCldaJ5HXcS6IAjPI485LCxd2Lp1
w2PbgO5sFutyaIsBYdsdOBlEz3edJFfy9HlPbdiIcXgf6i5/IPYMgOnrrkUkQnJD
X/aDbXUz3dD5PzaP+0h/2iSLmuBdArLqRS7NI/9YwB9dXnwOvSZXccIHVCo8w2Y8
ZMRQoqFwDcPufxAF558TM4NA7O6AfnK70cBxuKb7s6CCzw3EpUqgKz9QXU2sjZMv
YwBuKVbk930rs9oVhQXKv/LHPQ7hJRZPsQAkuzvnIkp/4cseIgKxjJwOB6ZINuzO
dwEHfNvVd8bYzx/G+Udvd6mHNhfNvtkwbHlNL/LI7D1itXzX1msO6HSKwjH9inen
2OsV51Avjy9kOQDJC7V1hyyBa15n5ZtoS6G857ZwKSNMqNa8Ikao4c5tZpByFmI4
xEbMZKRjdDn64X9hpxJUrf0jVfbQ0nThOvB+NcrZEHp29x0NUQ2gZDyUVI0Mbgrq
uJKgJNwyyogHGI+HNLg4/IRjjKSqM+y/3uSIN1MFMYdIWI+pI6SHcvjNX1ocb9LU
aPv5FUz6YnuC64qK276L1ls9LqPUduNwSoZzZY9k8ee5ZRnZemWLg2ADHSdj6vG/
X/CZQRCyVNPAhY1qkBwkhpp7QVkrRSiqbOeR1yPlE1C9iQ0Ge4BHxJguQECDZgJf
axFRyqiMUQu3cg41g9HuVX5sACPjj1z0SswS9ck+jTH+drtwcjQs9BrUz1RxkLkD
QbM3W5y+9CGFldVfR4FwVyTingTgVVTpn7v9Rvvtd0pHG3LYsGujV5nym9Pkg+cF
nNAninri1j21xSw4PJg6v0ZvV22B4N0qCQvPaGTqdyhXyNdK6OPSaVh0sK8U4ITe
+3gKDz1fY+9VF0CeS1P+7+3g1Hvb0Nv8Bcihj+jxIFxUTAqDwTKQYfP0iDEUNtos
Sq5/+8rQZovR96e883MclxACAQzKYgSTnCb94VYMxUiH5MPvKJ4vsozvsknqrmxE
iw3ERVGLtcHQcixZitbfGwItmWSa4ZVYnYEsKOWPxUjphByp1LFBqtI70Cj3h7h+
g+yE/hjRMEvBOW6nK8uoAGbZ7SWA1xiGSXlP5vj8/7ZzbmhzPdV08lNj/NQ5wWBC
zcO4YHlJnfYgpgbs5hHsFm4izKr8ly3bXCJqroKmkG7lTEoZBNql1igr371FQl5p
cbM22GfBgz6J98sJU5NWmT1QgctSZGPj7+oRsoD4lVEqWKMjESag7TmZSoLrzavw
sPDWV4t27tQuY5/rorm5VDRZJxECHIWnbE3xT4nDWdXsIjfk61guX4zNTrbL//KO
WPPu2GkFNb9/WQ+yA+KT3En8ecyJES9H/3ph2yWlWcilpoI5e9rJ1nEHkZAhaLtP
kEOONnoggBaa/TJVocyqMCcNgxw1giLNRAo/FnDIIc+wJCuoSKMX0FSp6E9PBs/A
b5MSigJfY1imadRUoAaieSlKFo0pqpk7UICUxGNDBcCKM37pBMpnuIuszPNRaQaI
NoYaLfw3euYPIZZroS06M0giIRJjyqbLS6xQegQWoUgWJn9YC8w7/gOy0gy+YxKZ
1t+lfL56vb+Ddj4A8fs/k0apoM7WKhoSbj/TVlZAzmzsfWoqQb31wkcVmuQn3mOz
7CtfhqjzeD9n1beJjxb5/E3ipvUvnn80kUuQ7cyJB9xxsIhle6thf5XfRPDNk7bA
7o47zo1pblh7OiTNtQII/4ioXNX7FUoLrisYGTPts5gdAOl4rfakvx58yVVo9oWi
74me3AmWwJAW/e5PWlsufjRPWaqUMUHzwR7G3wWV5yNhMF5LTxtciJ5fPlUla5kN
YIzQkjC2jI7niR0cPwiUrdYr5t9VfpR6mp9vA1uO1VwZwoiZCR5dDeOUJ4CGYc2S
7a4Eh/3dughJF21MZ/ZAm3jMomJoFKBXDeTAl0GRSMgffZfVG15R9AuDc6ets12t
72NMQAGdWtrcs6nC07tsLR6TrF94KSJEM5/d6sy+2mhsnBbODy6CNdw0IOzwl4RO
h6oXA0S0QpvOjAMk/+6uFFXJjJFDLKnm6VONG8HeQAHjsNHRRgIJphVsveB91HBZ
h4LDMQJ2waYsKlVMcrtzjv3xp4S5Xq89maUFEPpLJgJyZmjhONAI7Jsc5m2MbXFO
0yRpO3PzLMz1/b2I3Rb9y7t/x4TvWXD0HF7kBclsRFDpadnesK68FK1zl75bhmX3
QR++4UuqUDDJEQGs+QmpuM/4GRw2pzmpaRiwqLLGG0KU+FNArOh6FPa4o/OW3aI6
vA5dN4w+oBWL4KmHvyfvxpAfA0WbibHXR0kKn+OF0BkbzjwPN63Vhk0pHa0wCkLw
mNpiAnklVsq7MxxtLhjnHcvwclarWQvQc6E2/LeevGk8GfgNgHlSLCDqhTV/5Rg3
n78BD8xuoA5gN+SSmfuBZ/oC4z8KArdkxG/mi5LxNF8hfhY1Qqrz50ovYAZ/z/lw
w5sqaYKfNAu9deAm2aFeSjOAx8JTMuxoLSodNrkpLdPMvzucTu0GYqV7b5pbeUbQ
ZWukBiftB3CqMubfLismP69gwMWEPVbJ5aTEhdzrWklNy8jWOmwHEi1IGIRCyJOk
a57UD+1Yptlg+c2pVznq975C3un3+z1WhHflFsvKc9Clqs5IV849vLlH723t7qDR
4m/f3+mgFSHSynCbfem5JDrLWjnMMPKNPDsJjapuN5j0KdNjfc+MheqABlBJl/Td
z7V1suHk89yJ8tNZkBfZekzBNnR40Wk/1YXiHegudOPBhnxFXXdoKnyqTLQMuN5w
O0Zj/F4tfwD7zQVdgI+bd+1dRgWF+pAFyqeOUHZVwmuqlRIg6gGA5X8fbaK7/nLB
3joUl8xXlZXx+XM5l+lAbtASbKSmtdjzY/J3zJIdkIQbaM8QIoYIFZQnsnjQVXJR
a5pw0k4Sm3YtTtEngftV5ojtpD0McZzLsM0UQWpSiydw8CUKkkoErw40cJpL7/S+
mD1yAjQ1d62LS+cOBnKxs+M1ogYbChxHYI1CAnXGJxRBpkoAPlKoPd6PZ7+VnO2t
pI/GCl6sLtrxq7kxXcoO825cXKZGeyHlUMXWIpbw85BFwKjKqN/OoHo2t0Kbq8aY
HhCharH0Pnm2NBFOR2X872xvzQ0aFycuX+LfzzftmP8ExsKRf6xKb335DSkqkyB6
FaeTOkZWPvVKBG0qwag0Xy6J/ReEf2U4nktitvxVKJo5ns8lRwnHCjKHtd6/zpzJ
JhGkNRMxH+XyuUnQKL1p96i9206MeCXOaMtDpajCfkdp+IewllZXN4qfMznlH7tO
kRi2TMVQKT5wAe4qpXmu4QiNeiE2J5p4ARn2INNB9uh1LNbl4GMV8nWW8DVtR0s4
q8E/7UG1iL6GwbaYcFntskDBf6SHDL2Ut6REygsgq8wQEgTGifubQ7eVA4Ag4nlz
b+mM9dWrGMFsz027oLZ1W/tc5bha+vB57hlZXTVjf3NKymKB9rMuD3ef0E3kE4sX
I/c8lf2/ITFk8+gl8ix3Ta+Sh5BEY33LcXmqjpLOez2C9rOZp8GHt6F7YjCRNOXu
mzlZT3wSAVShnZMM3bYWo4nXWQ42O3lNGZUZUpL9mqMXXXcRctdbJh2Wl1DtD36+
7/+qlmvsr++8/B3zXLH0foqFgVmIV9yRIfrS5ABLgIai6CbpnRBBGGQRM7J0mqAA
ZvRlitjar7qlN80he8MAtdN3kJgCQ2l3LklqL3jZDL89A5p400EXPh6JBT9RxkIJ
OgZUtqqaDfAtPf5NOViIihTq1hcHYQj0bTV2sO4Pv1F7HJ4thvbW5iuwjFuRypFb
N4fdHTV7BMXszvCAAkUSn1Vauea+IVa2rpPbLGiKMVqI2mMeneZxqlDJTuZmMF06
o6aSiuR7/XcKb/DtxOKJEp8fE8jb2Py9cxsD52ho+oeJZ4a7t6LH+3Rw9foeXxWN
0cSjbk/kCoqve4+TKM8mckWFu7syjtEpRufUH+Db8gDDb6Hv0jiVdBt/mKd4RtG6
6zjzYwurs82F10WCyENOjJR3Tk5771YHmF34U5VAceuwBxy1dKoPjozELi0asUqw
URntQbYZg+yTGcUxTe8KAmIh0BUMEyNNKvZ55JeO4y3qIAIlqE6iLwo/KiO/L7Sk
thwMyxCx1Lk873Tg1kBY/cXvrabBEqsSh4BSUaEPGuKs9Dhl9Mew42biN2r2iGFc
mzYblNtWxyGm0YaMk5pwuQtUO91b8J5lSEc/4y72bzUYTjKI2QPyw/yXy+luYkEf
4LTsBmnEJR0DgKQyI4zj8cmKuztasf1Hyv3NfkzLKYJepQPGAv8vvRJnQB9jolQO
4/AZBByqAsfKlGhczjuFHxC2roq7lxdOTezqp5JaXXgWVDQ6ra9XdQk63HDw8wRw
/VR2EGRYnqc4en3MazI2piC39ECvggSyiAQMvGDanLeMs6RwbS84A0or2UElqy9w
N3N2tJ/9QQxKwlu3JSfyde5MgDz4P2eZj34WMq8aSp+iMhDctMNZj7AJSGkhP+Kr
XgGRxECBFsPhyRdbvSCHYYcim5u//nrINBk0lhXrsO+/6apWsVBUYN0Uk/a0/1VW
E1XDS9x7d95xD2+nyGc66br2+L+ob/zZlsSsxgUo6DXwinvFC3RtC633CB79qxpE
1ITN8uCD2Rw21PGl6m9ft015KQTkukm3AQ8S46jZRUcTk5j4Tf2ZCHx6RP+p1eqm
AMVCRiPs5T2jYlbGwfV6kZLKRhkvb2Y1c6fHgLDh6EPIpDUUg/5Tq0pF77eW24oY
7L5K7RuKxlsrQapy1IKCjg1f6AlqjDWT38ASBlEUXI5GiqVZournlVjm5RoHCD+d
e08hzobq6ewfCWHaCxLTuFNhWFqE+X97aEx3TX+NXJMHWxghHNFLpFgglx8Stp3k
4eGhSff6jLiMvsDUX2s4QmAwy3q9zMgKSn5jLTw6pR4qM1xwQ6URCnWvINoHT2gf
l5PHN2ZxkTiXlOO+u7BupV8utyT6496qyVSe2AXP9gHW94sR5DpTCgjDj8gDffg6
P/ton8zd3qqxWjToORVqHJCp7Z1La4uT8hknRXudP+/4Yz7guP9gYPc6n+PbzF/6
qUq6blnVQcAjZrxB/v7nHVIRhJh71/Tb3diXIrhdwR6q3FwQz9GfEoTUpFYUXFjD
S12fwE5C4dJKcqtn7Gfffy+zvhpCfQf7I//lJxUTYts4Lefxns0DODFRNXcZiDj3
cW8qUEw6ulea81Pnugn6OFiYPB/ei5hWfmhF81gVb8MxTxK/uZq9/t9Hz/JpHN6G
sYsow+5g9BAxtO0x61VdzUNdLqG1Yt9pA1RsoafIzB9yLqL+bydIrR0dYlAWK7bD
xk9CLCC7ZB+zeha6Qdv9/QBYifnuG7CDX+YRnGVCG88RBdyFAro5dh2qcw/ZsOGX
Dd9vRBOkrtj8GdrqXJIwpMijugR98h+Jcje7t/f1rwjgF4mlkYyLtBXPSjUBFlxW
vMvl/aKHxnfRePB3kgn0yY6dj6I3fI2/igQVWY6/CqPHtjS8ErjII73sKNBmcEOn
a4AoRtPSGLorjrOUbSAkEa+yvObcS/TCphqertqfsWQ6nzFnn+ClXixk+nkWu2WT
RjWaV218RfM92+q6J0xhsfcAtonzzAc4pqEkxAMjx+z1n2lgRVSOXLRwb2qk6hs1
3iVBvKHNcmrT8+C6Mpj0vCWS4RkY9Q7onJ1l9ivAYsXXOCeNuXk2yOjKdHFIU3xj
TVZXqP9b5i2zW2UqhiRnLPWTKWkpInZ7gUXKiWaCCAaVrYQfZKCJdwonj4gYDvj+
QwTdOP8sAl2eAP/QMsVlSwfI7fxdu6D8HG1Bi7rcEKJMIffKKKE4MqAtu9oHBYGy
GtaxJ36FOMcY/c0SdXAgTMhe1/EqrvNJfRl07YFZvRfuPxVaV3iNIsabxPXmM/B2
W2DBh4FqMvtVPwNlBrjuXgxKeAMUKg83Lna16gWMqhtuBfmLrPD+1Dp3e6uZp33k
a4eQOuVUzcCtvkrR/an9xddkIb+DB9Uos9QwI1Uwe2m+gIp98NZx1bz/VTS89EGg
NBgG1SM2ijtplW1TBoSgPmbYSGRmBzu7Oo+a8gHqlLU5tf+NosVWr9l4yCEtJ7GU
/z5fNixyA5QoxxSGyqBuNT6R6d6gx5zMNZuKGqtXl6aHFS2k3Z+U1eqVh7hWmnQo
ZjMQvfKEk4pRt/MN/5ogUu/mmEbihMFfUsGO0Xm53t4UVB6YKPZv5J6cLQ4wdMQm
CLc0T3BNbiJ6fMPCg/yM0PyHkfdXobXnMbsfzRQ522yEzH2sHupsQXfj2007GM1j
axx2kO3qguil6WIl2jykPVHrYzBjDfqJO1VYZDjLicLDMJ8/X8+DUun4DO9INGrZ
9l11OKSKPgMgcCunzz7cAK/ZrOOxbLodBZloyMUq5WyxSogV4uuDAup8KjPqqoNz
J8jDTIuODD6OqL+7W7xGyAkC9BOr0jMKya7LwD+nfpGhsKUjszoUwpQ6eJ5wrbfM
2Fp+Nm/f1XaqQ68oNjMuWOuJcbEhALlkQC5qMRyeu/vQKILcdFSWXsBtYjqKC2WO
2GPGNa2HNXehCcCF9kesEhhNPXU3q9ZJl9gm8RbNKkj1fVktxJI2W7sJCi/EXXiV
9mYxM4nigjFPOLnJ04pJqnCPVnvi0dPotRVyOa1/J/QVlQkH+W30hXC9S7MxeIX3
dVK49h2ETJqaDHvucujFZYh65ma+GIfak1fhzAyffJfZQNAO/uAxVDgN+a8sBQHI
rTPRqZp9fU9L/yXnjgGy46zndDI50c4kHCCUnLLD+ObIiKy9kuQsT1lDR2iRuTBB
KlmKoQQbDFn7in6gc+e+NN5c3aKthUrUIlsTQrnA7CMGdK7uTU2v+HETWirNOgaV
MKVhUvgrsfG3DJxBNfK+96zDeCsZCFeE9lzqt2OQp2SFndJhzySAZQHaZHcxoCt6
DRu+USKBXpLoU55D7AqiSW1yh7YCxVITnCffLRi7auSTVTzEvIIM2/JGRbEzvV6i
CYSusYAcxKtKICKhd/8NqmszgUNmjbpWKsu3q5uRqZxaTb7D42xtpIwnrDFGVc/1
ciUXezPpl43kvVfiKcdoehc0TAqo6w/iXXGx/SirXvr16EvNFbS8DuI3uF2Cj0Us
k+2DdH7ZFqwFIoytDG2nE0qIJ3kt4cNBIqr7sGDVo9ICiUIxdE3/ac+yZtrxpKeW
C64RzS3w0JenVNnRlV6dkWpfS9ulYcCDYgvhOQTGIZuyqb7s1pwcHf2EAojWjaa6
0/wptiNNqg5mQIxjl4YuW/LurWxOjuQ4vyzhpNB0HoynQrmyIBS7KIERwiuE9hCv
a7/RiFrWxDineWz9eH+e4lQC3qdo8qsCI+t7OeoYbfCxWJN7mTcjrBUh8w/XiM9D
28u2/GegjoSWjL4olNHeQ1xiXkXMqKucvj1leqZnDdQ45ByUxzABRefLVGZztYBv
D9x8tDtl19pix0qJunQ+epd0MECdGghxCaSELB2YwMsn3DCZyBFrk2+FoPK5h18g
mIUx91FlloJcC8o/olGAHs9/btd7/nLMqasp0Tj4fXjDthXi7SuKIQbeLBeKdcdZ
jWAq7RXu6YO/DayU/6XoaSt7NfUXnFb/X2osajN84ORk+Ej2lXY1jIC4C1pC3UY8
CSWYK6lZ+sDVNKKtSzkK/AZNR6W/CoUfBsTBi7eBWnJf4r7sm/UOP6h8D5AFOt6a
vqp5gWX2SvK5dmiUIRwRvIKrNgZpRrSow2tgWbTiTm3Uz6QGdjuq9mYW40+mrVmO
W6EncAT1K3gP/2nG6ITHsF8RWQ1/oZbVLkqnjKmYK8cC0bQ+ofUH+M+2W+/IJiuJ
guN87hOwaecrHyZFX/2L6amZdhYJEFZTZ7LcQjW6pNg9849kHxDo88eZIsrRlDnp
rJUYj7asq6xZ5WpFpKb95a7w0U80HQ3ipkZVQ/NC84oK3QzftbFGts0i+ibw16UF
k7z6cEqxi/M1TIoK5Ll/DZQO8irvtiY2AoOv33bdWlJGYi9Mx0c36KhAevMk6Nhz
duhHq7IU0IGxTJRmT/he0HCSQ/C5mQ4esMPK2vWWu+cn3vzOtSI60nydOPl62qb5
QylZ4kponcdLDCaXmvQefhypVq6whHepCIVYcSMGSxuysBYzqEWO+Q2rGemxFcrp
kQrx7Q4G6TZAkxeRTWveCeyVoC2pSEats/cGysITs7CQBA3CIkJ4BMufpvMyk5X7
9GktptlRrsGaKz2UdixKLArsDFuOunEc5nj7P5e70xZ9olCM9N4wGYQGUCHkFlbT
1I5FrC6NFM2xj77X6Qc0mJAN+LZMu7OUUog8650JyM9++fLGntQZXNzptWVOGvQb
qamHkJoRH4dPRnahclQZanJQlvh44lRWJqFe/idn2654fIC0ON9YRJVTbAlEOWyd
mKXUb0kP13yq2t5xxM564EnmE2bdfNwNCYIZqEJ/Np/tGUT0kcUhAJqDjYhbwupf
fqpxoG1zskMV5nm6fZLU6JsvgV2h61gJrPJZC1E01Sxt0XQ5778mOy3Ys1N8LTcc
v1UuhEP2jcwpuYxahBQA9fZqztMK46/Bgkvr9hcHsgh6TQxkBfaTRSqxka2VBlsF
BXCmFEiiDkRJGC2pz+7jMIRp9O2+Hz8oGAH629jfjzIokqw44b8CMpMzDZTMov5x
TGw7CguiucOZEGwYfkyO2jUj1XligBfCFDM0JkWlycaETVLZBFRcopAE/KNugIin
stsZZxTPE4VlGVGSdch2uL461u83OztnW1Ev2dX9zgj0h1v81HSXrXdJ/O8d8Lea
Tthz8jBoIYdMK1MLmqRDEEMLiaMNV09EqKKkKSh16u7G/bLukITcZhf6/erTiXl8
W3Y1ja8PmDXq6TatAFJ/Mq2lAdcAkfCdET+dgr69oMLULSR4yYsECi+FNu6oGlJs
FDYeOhiHdpFaJgsAiicSp3fobHtyiFLftt1g7RykZ4kKlTeyIg77KQxyNBhN8coV
ebcGmcUtD9y7fLlAPqkE1PoyEgGuldgbZaUkT0fIVEJUIARnPXwWg6zazBQaCozt
0XUIv/RQfmCw5vtMyUW+pTGSL/L6Oh3/sk4svqvAgTFD9SaBEoOtRavjSO2egPty
7PJUaE8AuQFD8zXsuOGKQ7FuD6zAtNgjgo/4eIWnTgVZAdCw+CWzwlzNfa4F/LQ4
pwirZuQcHBYbw1n0M7J+YLDMqSSn7xS9au+yh2QnTep1taEU/MfqsMA86ZoghOlH
LjC3rfd+ojf8jOWu96gaaJ0qhX00MenVrB6H9kbcp9zeM7nLoXbOZAijKmdwUGQm
VvAwjohD/u/scDXZswcGO8lrysDsWpsdieGDcddN+Qguc0pcy2T6S+CFWRXqJyOp
sURKpnyVG89JPTiYMerN7NK0Ia/wXD8NfyNxYGzAWgHXSuzqsnMCJD0GuiWcY4u/
eb4BBwQg45tTD2pIihhH4X9uIrTG2E/hX8uYnU6HgmFgKP/yJ8IrXo7K3OIBMFyr
0IAnUTSLgODLKo6ODim8M34m1eGMd0yIwRCGCONSoXH5UlEkk+tUBgGZMj4oH4yp
HSmPoepA3xCJcDE8BQcUXsw26z7Af7K2g9rxm+VXAjqPFBeCPNvF2XqyqJfinS31
D5CyD34uDc2aeSMWfLuXfV7/4c1t07ghR1Uy5J4xCUIG8PEG9GOGhtQ6Mw8HWkr3
6cii3ZGADXi6SCKywtQM7HqqWLT4fnqrWFU1QO8H9smfbKqKbEqbOB6yzlyQdAf2
csayfGxCQYNiq1KXWvPmPMLT9gdDLRFLdywN2bgd+W3X/d+1lmB1xr85dF81pvPj
vGN5e6vh4A5KRAs6Bon2jzkd6ks2NNLa3nX1nKaCmlq6H78QUxdqgajBYsUu5XBR
ZI/RpA6NrcNIykThTMLi/8DTbUqpHoDOtSaRhZWqN2JWFoakNvo5Y2bng85rWs/B
4OSJR+GzmyJkgXprlUr9WYsEM6bBXxe8f1xyst+fXf8mqqZKWpmCHLFRpTF28XKD
IcZnXmGu82MLl1s9EG2MpHfXoCvg+QtAq+bmzcuFy0SvhQfj/FqkNo1ziaiU4cvM
0Vsgv/q9X9wAtse9M9lgqrtgPWk7oHZalWOXj0rae5d+44Jtm0O0mU/mIsqSUDC5
1LTh1l4wjNiitW3di0sIzmDoRhrpX0ogipcZPBlNPxvVLsfDwalvyk9c2JtLKAK3
ZbqIbkLQy18ZvcvFr+F/XN2q7yB14NzLMP385B5U4VoBHXlfE2yOBa30HsHlwhtC
P20H0/7YcZ6qO8o6FtWPmOF/JMGCFYYyPn61sHK/psNnotdrPly21Ms9vYG8ghB0
l4xmLcWKslYvXeQegx/QQqHJwB8DpWQJxNQI+dOkl3sTznzKMY8UPwxPdldJ2b/2
SD04RE7tmFHFyMy2xWo5LZejTHVFUGqA7kGKSko0qhjJxnyk9Ie4fLL075s+7hV+
DpQDyq2nDB4BJC/LE76ITf5YSYRq8i3mm6Dr3b/OzKKPqPdG3sVn4ftLjk/ANxj1
UTbIMOC99rN9gRjFoswrHV/CeZQGKlXjkh4FEyfWnx2BBeHMizotwGcAghrziBY+
R9DZ7Ov0xsfCopG0sEIfR7nher19+r+YVa1sgayJxFRJzC5WNhLPHHI1nBa1lByu
UhRqcXOqXPX8jgVmR2uSZ2JN3jO/jFu2MWOtvMExzfGPSAJf2ifdoqifMAjAuFc2
OdJvnTqRbUD/xjumyQQxCKrAzNu6X1497kneQv+flGZ13UHU+H+8nf6r/daL3/Un
EB1emluuMvWLkQAzsIzAW1VXle96VxRYqc/ckO2wNMClFm/C7bYIowhCTFhNLhpP
Or9v8HcjkKEvDkg/qNsqMl4B1CnQe9ecb+GFyYxG4K2LRt6Kg4yJqty4KxNXQjIw
TZgEwN5/EX5XBNzRFFaktt38HnymMJOrybzDGzjf+bGW/pXYAWbu85xNeJM0Wabs
1xYMcjFI700aRFdQLsj75ipIf2XH5QtOh46SshYc9Hbe/WSFBHoUXnUjdijRskT+
vn2pTbe9Ut6fnWvtV7rlG8NEAGLt1DAPG3O4crc3spgosOu0qzQ3nTAx+nyrHv1a
BuW/4UWdiNAIYAIyTqMYNnz0u/WMtaTFvaz6FJmuXrmNeShL5Bo9sstFgI4+sQrl
IuFJVTsjY3uttsmL2gRC0MJjn4ZTUBJArmA5r9GOlH2HqPMP39ic2x5XdfQawGHF
ODcC/XYrSpHdZpxfZV2/Qqq9QL4brEvmtqzaOmOX23xAQnrep1TSE+8Ozic8vJN0
6bmR2USLawXFooOpYpOrgT6TQuhKJh/DVlmN8QXXSbF2+NPqF6Y0WgqsKzGpfYlH
LcBRkOgok64bDMTJu1JJ61ZPiYurpV4zpe44JCnO6QU/Pbg4H29g96oI1I1QQFSA
3bj5jGOxKxyl1hytQDgDnKU2lgX2xHPI2xnl4Zgu1hFUezK+RLUnXHNiiOjKLXda
pvo4H6Tmbm2GEwKJh4aGJ6rFcdefiPP+8T2Uk+CBKhhO+8DXAc/imIxgjml/i32p
YmI+N9p8c1+TdA5fJcbv5qTL0dgE1zbMeUqNVaoDyIQfe2DVUjTWuCILj1ZKXiFs
XIwkgyfGB1vg72vIPxKcxrTLQcrg4JE6nu+8zAlVGrSZ1i3M0oPxUT2O8cx8STzb
H0/XpWR3LxqNxdQVdl6vsgW7lcnZfM/zCRE5SYevDgwmKiifmGtnYFdkSxt72OdS
C4PE/gk+OtLVJWqPQ5UJSs4vS/c/pctQ2nPzXRbKNM9iqY8a/70qupEoStIZ0HPr
+uwCLgv0K/lwlNq8m1LJmTDzHlmD4BsPyoiZTXgyq6pF5Ix88SIJqUYC62MiL0Jc
IsfIMxJO009NivNdEO1LyW+4O64yw/vgYxUZ6sp4n6obtr2ykb9qsz4uU/4xXjMI
dFcOR9VyauuXSNY/yEX4FmcvzasZ/aKsLtKPZa2agCiXlvCTpdZYOvwhn8VXd9jM
anSDEfEcA4GaWkpF13i52bDwIXtv5XtKbm3/9+ulxaFP/Heh+Z5WHwUUJ8T7LJ9w
jqhLXzlItDPEUAeFssg43mYVzt0V6H2qe/L2ivUuQuurZOa6WBheVTuraIoF6R3K
xCVyyFWmPIz6kN5B6nOZNxOhgklKfRr3gnICylNqcWFJNrsgdyiiOM5z8uXWoCk2
QmobwIjure/pFlFvZsbVWVlPIkBq8007U8+zt/A4MGlaVzwSz4J6U+LDG4YcBr1d
IDRgpNH8LfjrVTSpZOPImHZMTVpeLnlCCLtfmlht2wwtwP9PK7STD8Jb4GY0/+md
Iy9zv5RxtKGWicQBQ7Oa6Xc4FGs0CcrWRkVH+68LJLQqZsYzHOOia4On6maIe3HV
/UFo4wKiiIlbdWGBdAsCWNAEYagZSF5VPZK0zWUrSZzY+Z1G/dIA3AIck7RZ60z9
zV6p82/y8bRrjQK004RtrJIGeWy0B8GfWx14eFdINSAkCWNZ6Sj+yJsKVFigiCuo
BPJZQ5jEa3/UI/yZk8AEuXVhO7KEBot1Ez9OHkkSuUJSjRY3tVsLS8efxGsz04px
fkb7Fupwti+u8+bH9qhfapPafmoMQyyzZardp1SDftd8jUZrQV3YHJKrEioXBC49
3FuoZchin95f+7j1PjrvIIzXMH+huVAr/fksafxSLrH8cBIxzhl6s7Jit0Wd+6D1
Cnb5g3RqSkTAzOBd0s1Bbccvsw3HI9KItG13l+RMU3eJ76iSDKP1quUK3G7VYs7E
xGryIeNx2ksr2IofbaMG3dV7iOfE7INKXaCNmx9nxvZam88ob7HDDrTi9Fe1UTM2
CJnpH5RUayueKAwG0JdEsSpMKuuvv/ztFI6eMdzcQc7dwRGrJQkVXNYF1ji3ykwh
jjySODFu2YiYI0mk+3XX9UFzSryvZ9hXNKJfcsxO5c/0OiSIEYdmbflXGRG9elT7
YMO6Hiwm7Rf663R5tXq8RdGTuBiVZTEURN3dStVc3RlrtiSvCbTCavCWK21N7NH9
uDLO9CiWrbWDbZDjvh50nrPsphFYae2A7cR2h3vEvQxAb+lkvS/2mmfh/v4Wjcen
mWc9TCA1xmALndHh+aUVNaMeFnWQ1G1pkP1Yt8aQx4ahcWVnFlbhT69LK7GHZv8B
hrRvYTIhCCAZDB3gf93Ke6O1fMV/WK88huJ9Eu2INKwVW+YZQZv/ZLOX3Ic0IoZg
JPdbjRGRQUCq1/kH/MisG3XTSI/eJkEBmxIyUnDUBQ2N/qpYbx6W57YWHRM/gco+
5LzWisL8eTPLoxfbh7KUHmv64fNxJTOQ9Ak23cq5oJL36SQ9nOK2VAOk/FVXkVa9
4TcgH5HM4AkEki9ohPdUxFUDSFLnjUFVOiTO6W+SeKRrjnn0OQLCCP9qgzNjtSsV
tzc+lXB75xHya4NaxlVVs9Bp2Wrk5SDsvM8FiQen3DIITEgV3YB7qI5ciRNaiEwL
4fGtKQ1FfjLekgCFWFFi0JdVMKKxQwNKs3Fw23Hina5b6k3tqMe6Gis8nWKq815I
yDlhFv9YkLEV+VW7lRzq413/b1L2HnAELwrmv1LR6ZIT8SABC8yqpyICncC0jZaK
doA5hBEvMxZaD1BTI8F9c4TIfHTH9hGBkH5J4HxYgYi8ajq12+Kgu6UwZC7QHZge
qDHKWemA+iNJNOoQODqwNyaFVIeez7xuC4ghhyJ7ZlB4pAV40DF5lJDZWcnFuWGa
Q8S4nABfFBsx7D+1vkm4CE5Y8wCw16FBFvf8GKq3e+fE/z3VJXUXCH462CLSNYBr
uk0AxlQSqjoQc5mxYfaLVMGgTPbacqNMCJ31Vv8kXR3odmCTK3yotD5w1b5sbyo/
oMaPR1h20zn+XS9jFEKMYOjLms94q4rjXyjZ33OfS7/KWZm9JnTwiAEG2tGcgoZS
qAQ3eaIE48pWn8tHw0JyFeH9Wwi+N5rkfhuVE7HFSjzVSGkmwK0E4Rm5Jl5IEKKJ
QfX5jZCHWbL8/OtPlx8oD9TlssFm1B0jE4qscGNIctW4xOQ40KbDsy5gGdrjkNec
q3bBZew5cfT8w6I21IKdWP7GtKfePr7aR+NnKTs3Zdu67NHgWL3kjToFm5JCy+uh
CMszzgLnxGY7geJjy9sUaNCUjjYYaq0csbkbnAlT7cqCropiPcJ4Pm5lRmLWMWRH
IjkgMoOo/EXmKAhaqJaG1rBC4NEJ6acV9x68l0JyI27REhCCYlYRfP8tWlbbTQl3
K5awQideopUVBYaLHKdfJA6fPi3McoJO9NckimlSuL5UJGXRUDvdWaCaIC4NNd+0
VhRIxYcRZOb4lTkX4qwLkHft7o0iujE6kc/7vboureKw1E6CmcugJnp38ZPgORA3
blEKI/YMDX83Dsl0VA9pEx2HOyh8OVdSZTFPRVX1pHqSgNGOAFKdxTevnNLrW5hm
097BP5FF8DHpfSLuvVOHtEovyUBpP2T8qr2DyVqhRLH5hQXrJ289oMtiqul7XPiA
9a8LyFkQa30/wkvs8rKoafsOOrklnqvXy+JuoSxo6QeERNYeRCCWONmVvcjTK3a0
d8T2npoKx7SLsfXRG9rLQ038Qtb7WmtslyYzPc9kHhFsHT7B+Os7F6HAVvMES/qU
b2+OfYlbcqF70fecddSHjsdxbwvx/5LvX6mn/0oAMTrABIwEifI+qIOgDH2SI12K
EdhUccuxVkyjt2Fzf33N5c0PcQf0JmL5A/2n11Fdms7GoNvWEBI3SoTJ9DjyHi7V
zdEfQbhi1qarZ17lyuAI5rQAeQ7n19xp63Mzzuwkujuuvn+XfLJwze6R3rPkK6aC
f6gIZg1JTQ2WQKJBAjn8ROocLWFjAx1NVStRcU4FmrdOjL6jIRbg51G0dHsNMoaC
Ht6vf1i0hIUUd/OSmCsLXb7ZizD7aBJQQnmafb3fQ05BadidSkzQNMUqp6GvA17f
W45k3dWmN+Hc8UJaRuceKC1sflMxJ7lqLaQg/fmsIMOfwdCdckYvGnFSQinQzL0j
LmX8sWPCqv8kRlt1HaZQrVJv1aLUNxWlJsjnQUFv/Nv6c43qF16iqrdtE6eYFimv
yUDbN3eZMDGUql+5l88MpEW6D6bhflBYZOrKklivZmmc/Ce5Jnz8UDf3+wfNqPeR
/nqg66NHZxuG+xrt6OOeTHphIsn/u2X/nBIf9a4cSfvFSBrdLNWi3J23fv8AG9qR
hUEw+pYe2HsQXQW2ZOzdEp1103SYD7gkOGMlJ89xsEEug1ArP3uK2fPwu2SMPj3v
V1CLmnlQ/FJ8Neus0wIo2AYTztiO7wjM2z7lKii80rHvCOfJLweB00uCVMzhayGQ
dQ0FNxvooAmoiEShh+x0MzbBC7g5lbmOTmDsYACSN6Za27vwMFPLl7HDwj2n/ByO
uvHGkqOPMJmDQaYJS0rFqLyHHQ7C2swi2lzAx7cIgIzJNa8JSSjy9CCbLqTrse+t
fvyt2+p3HOrcJiqO6NKJjh9f263j9g5i5W2xcJXqd4HEGC4feo03aUdu+fn2i4VA
YB8axIou0gA8pTevHm1geUn9wSDiklbhEKcF5gSp2cuwK0bkZ2KkbJIwwJHaCWn3
1OQ9rBLoqdixxhy89Ey6yyh95UOwOUUyjDErqqprfjBpcNQW88plH46t5k3Vdfbo
Cpwe005iTtc1PJCDQyXkHmaCMesa0b0jjIUj3SE4VsM/U9L3DSXFb4sDz4+JQqvZ
fl+/XmpNAQ0RSUQTe7aAbvHQLNDtNX7gYhrpRPj1jv4+VEBBhiX8L1a0nghg4igL
EzQyaHk9M8UUvwYQqivkvUTAJ80glZ8Bksa2G5yg/KVHmTn0rzGHUVteZc7s348b
LWI7z5PFkpsxQk3QthvVjV9LkHBOWjrqR5HUHkqaISEPyUjQl7P0bcgiQhwRR9Sx
gOzyaARrDkwlH71ubKXgqRYrvraWNNPmCj/exc1tdYaOveFKa2M/LdgDWfq6wMaP
6hhVMQRjRdbxJaNk2QrehIb9DyO5Tj83w2HYKwI/IVf4TQmMrF7RahEmG3vcC100
5D44WSe5np+z6rFsPfPd+NuNNSlblEC//MWrUdYYMQ4WkkzW0+N0YSgL3vQQb3Kr
1nBBimPg7IyvESU2COtXJsPy3W3Zy9/Zkrf96OD2EQadYdNnFHy1Dj9N5qLsnkOW
4MVwF/6GbJywDwZtVNboqRObUN3qmqUH52M4YcE61NIWEDtUIL1SjuDt0ezk/nbX
QN2GKgX0efWJD+Yg5UGVASvXprP+PcRM4xTxDwe/kP4pdAHM+s/7cwpxcMJk8Tdu
hRiRSWaksKnfYLV7F+ySfl9f+lR4bTI4fWvik6/spL5xa4ducyy8PplxBi4CxBpb
bTHsaEmrk5SMqDchtfJHOyG7wJTYLL2a8JpEwtXdvs/tnaiqZZ2iZBD8Klegsf51
Gjzx2ITXZHLH2uoMW7f15yOirfvmxWG/lTUjFNz+sTeI8wHHaV1CRT8PeMD6Wnyk
fkVlFQbqYghyK0rGIW49VkudMIQHFw1TSV/lbP8vp1fxV4bfmREn3Xyt71BPTgAM
2888FFMUX9PqJ+lNTC9xAdUv/yqbPrUhIE91qc8AROnTsW0LcE/xMeXlHnwqpJg2
oiV4y6umU5U0FdD7oyeZSvfbtkmNcLx3keAPUKkarpGS2yZY5mLP2tIXOzMEtHsv
v2v51odeYtU2+SQB+QiH076PSysx0fc7s6rt/BB7F4/yF/p4lD+Kus9ibvrsYpAE
ySCX3Bnzkds57Qs8BDOcdtGns7+GC5JA83XY+s3A33nE4vp1yhkQmGWUit4tbD3d
y4z1kbGrZaW1P6X/0zh4zq7/GZZ60Ca9lLQuzKx6biazUDuagSu6voQe67r8jsyY
auBsnWgVpNpQ2TBCmMDX8CfJne1XIuN+GhjwvuwBdwbnpfo06J6BFAssQ03RjNb3
fi8yeA66Jya+lp1Fqo7Va/LTWLydyt4kbc5iix/wxhVRJVaeHX1pWcMYqT34X28e
eRqOvjEDdmHz5gAJ/ZoD3QCJJiSUeBuTY0JoFamyfbg0+GiyTj5ClOi08m/LsISo
LWquzdegScNkXS81puCxSoRrxv5p30BfpbK72nC35bd3OL4y9hnKoeCE0cZw/eHb
HfjDSVoSVaFZ7hITkk2dCcYdIK/7eiX6eNsaVuBKHisJzL5XEBPkAvipMYbx8abf
+G5fTrMWrPbItQMmuk6vzLVYhpZ7SD3IDV61Obn70B8z1ZR/inSP9qJPVN2vt4S7
w97J+txpg0RERezzyMODKcmmtlz/iBXzldK1SlLE6qtCrBIsFaIeQMyV1UKxX9no
UqDcNoWxlzyWivnkPjxdCD+5lv9N5PTxerYSrVHd+ioDX4MtWfHj1z7xFhhtEbHz
rvLP6mDy+s7jdV4L3cXwZqPR+ivB7akZ9ujrYc4FbuxvHN4Hxhpl634hv5MEq8Xe
IAgGTC0CUtFM9TTwtpIoFpdG6O6wqe7bWVZqHo1Iw/LMd/y7Od9khseldeOSdzxd
J9Wyxmoi5l2A27VLaRo0QuAeaIvoKxip95T+GHr6G9mCaKmsjumJ57kBzWXALr9K
n+ziJqTl5A08nCBT1/Ic1uahzo3vMtyaO/2wzFbHErv/T9XWVkBA7PwshzhC6LYp
fBuZeEfQRGN80kSdrckmSbu2EMmr9vKU7TFK6AEav0tfDnVFZCRS685pXR/WDlms
UGeQ8OwF2+KW4hb9SNj8V+bYhoSv34iOeF88WE3NNoCFnvw31E8qRjh3yrO+7Dku
MX4giC6AIJezasw5w+FdvSSM+51VGPbTvGam0yqv5bhjLzRVUGRlsR2SMbQpRe7h
MIJubjghAW8b8/hBBxq73NQV5xdHj8mOvXs4x7+pDIdrgKweCUr9gB9A8t51OejU
zcvP7jh0aePdLqlw+aaNWTfUuHTKFM0+nJojHfpP9Q6yebh0cmN79rWVpilnDTvI
osEZQmni5eTBAHyXYPfhXm1T7eVc76BOK8mF8socyv0diXDVIvQ47wtcrO/pUITQ
vOKwIHaBXcWJhnhqBSVL5aznDhba3r9Uyoq5Qimhey+7AFKoOI5GmM9xPbUds81P
GVXylJBQp527YSte9+2/FkbFZTRBw1E7Dbech24A/rU+7kKFZRnY4H/v66oECrkT
xSXg3RYFDdkgv0f5cr0LCS+u95F38JgcP/p5bNc875kkVW3+VS9h/hy7+WfnEKX5
TRWz6oY0ecaNjIkxfAP5cLfC30w+Qqt2v+G8Bm2o1d5vNs1kBbWilbF4DX3iLZT3
u0jxGuj/0aNfDEV7YeRZzxxqGJs9O+jVwsBldKaHFxgHQPvBztf6tgCHJ5itYP8m
Za57B/geBQ9pB9yhVWuiPXwpbzRMQzidCBVE45jVEokXMDXn9clV5svIEFyP7jSB
Mh3fzqWP/gJ9MQ2iBTXYrpXhOQopJ6eHmHdCSSGEC8+VnHijMtQzIyWipkoZ+pqn
TzcUQfXtVGILXPjydj/ruR4NGaSeSnly3mx0vXzY+evBwVUPrkxJVKiBN+ebHlvk
8AOcCmPPPWSdcgQ75tNuciPxwffFq2iAFCTulyYG6OkI7//SmKQSitzqWpMQxeYc
vtz0bqWdG+tgBHEcjijxhYukggX2t2UuziazQAV/m8Q0ZlWpMiMXhymMNIakoOZF
CW4GuCG3a8sqOH1fUM5hPNEQvqLK5xgc1UYozQ4PnsNTAiY8QfjpMIrRdk6IDz8V
FE0LDxZwIu1A6PhS9jiNYDrBLptLabCGp0p/NWhMQw9/byEVi5NE6iOnnFd4K4MP
xlZZRo4r+SWge9LLA/V+0zFajIp9D18aisuQeLh9wBAmyiYHvN9+D82bjlHxrodd
rp1qw/vNtI3O/JXjHQDAuLbPsEF2NPp8/g0imSb9Cy7FUsgxsAnrDbL1xEdBR3Dd
1b/LLdbeXD/p80MQslkzdvb+Eic40ge20GwRKgPmc2jIcZE4lem45qVz8Tgqca9j
WP5XhuNsSu9P5dBR2BLecZqhQknS3JdL2vkHNrpQfv4cNbczI5On3BfggWtrrFsn
zxvuQWdXQ35/lltYfm5sDvuEJIE6BwJ0MNtntanPtP9qmnmJu92GwUqH1U+0/b7z
xp/GJO/qyu0MkYLh1AAlnjx6Edvf/RtHuIXxcvCZXRZRaSLMmfBC5xl/rPU3q7oW
yTY7BHxswd4nQw+HUJP3LpkZkME0H7CvXCknTW3OkfDf7bPyL8MpSAodKQthIUKa
RE/Unjh7a7Y9WktZu43YwBa6j/vhc6jMG3bCBEI1m373WZ5sI65kjFuWXZZ5ZhUe
1kQ+v4hJU65xGlFs9vlmke0JbxfnxauvJqH+vYxa/d4pfzYThimUUWn0/rW6EbrB
W53VsyKjn0Utyadc63p5xsyRrh8GjF/rFIOT4sCmbzet74u2ezwPC7IxtzrcYeLD
qgOhNvU8oBeosyax3bzzPdcs5ATjAX2LmRpXCfdDh/rmxDQ5uIbx05o9NtbEd7jl
1zNosi/L8xA3GkzLbSOne/WF+P/0+2vei3a2zS79mbGoazDw+4j2RkZ5l+s1Nqll
On+dgNHZz/5p4RwEBXVxWzsJ5wrW78UQq0lgohMv5gBq2EY7/6o51GNJtPHuRxAF
RsWuUgAF00rIRC56BgyNlOnkiUrpaRxhpBJ9O5Lzyjk5Ju2cApwTH7ukaG61pfOI
8Ww4QRwD4mxYniVKVu+AjVnAacoiG4UzaOX1ONsaWpNfeqTRXUhWoTd7N7aKB2Fh
jVcxb2UBDz1fSfe5zxe+Qh6YBfrx+vRyTiiGYB3nWp+KtEj2JYXLU34+trwHiqrk
lvknxQSnuuxMpD9/v+xRiPRqZyvdRdiV9TkFexh4pe2TzWJMOqCUlB9iEvCUzJs8
gcPKTwUqYFJKerLSuWQHvRHr+ACFzI+VdlWaEe+BY1nbjqjiFjdHnf47AEiU8lk5
V1QtnQmS+dRGWtvq0D6xYlZ3aaoy6RKSjZ1B1fKYu/fej86AHnKPEiuWoL1s9MpG
pA0ruO8bCh6zP2Q5PvtpCD4BtHL31KUSFsIi7qVkkk0HG0Kk3gN+ZcfQoKyPHUHN
gD4fwLOP2IuNzc5vvyrS0lOmi/xOFkhyuXm3e12yfOXRwBRD543RsqrC3o8DCeKE
I8RyoAoX2geOvNk/m6dSUpp73dA3c5MJWhTi02yNMN+ju57LXfLT/D6Z9eap2uIo
z6MWRG3nBfo6vZfEi3uPSCyyvXY8bpWH5Ga+ctQ1BSfqRN3s6FgGqbtltSnRBwUd
s+EfLqHhd3IehHKSUbGFuK8jopc+46ig7WOMdMPFqeVQqEHlsbQz8qiz8A9Wj3P/
BFg5pknByA/njI0WTQDuz4Y/CWtmdiltrwFdNBI9ZtchP+Z1vkLbEBOhXIZEilPt
nTQjLYa3rpgkeOQiG+5olTT0I+9jE0Xc546teUoHS5Q/P+gCrMO61I3IRPJM4b8t
UX+tieLZd2TYZK8d+FXNJ6SJJ1y+/ZH2Dj0cMNEKLvIiojMs2GpOF6QHa8L/Ighi
h5vKnQRdVxLJ6apBJA4iW7Bjug4Ffg8LsDMZckdm1jtUU30P4wwUn5bV51y34tr2
CiwvTWYaD5tH1NZOzrmsLY+wQGjBcqmjl8xV0N7I/Au3l+dGX+30kvRfm0Tcclc3
IE5/7gNtK0s4/moKQSoDED7KV/qftigI10yLKHc4xbpEELknvZahBSHfk6NpU330
Ln4lp8w2uRl8w2arSeiv4A/OA+7lvdmKt2bzFkajyI4DNmVt9xCTpn2RAyhh0E35
n7LCTHokGfIRG3b8cCI0D8l8URf528oSFRePJy9DImQpOUjOfKdfju68rpOuZK0D
WYcvJtnvc8vHnSY1y+MU/gDtllRM58buTaZhgXPF2InuEEKWgQfpqEbfrYMDaBS1
p1XEoOV8C9cFuW7585fRu2DbkX/tXmKU6aYJVP7PIZeu95HFTV7EV6Pj6//3Eb/i
1qy++DPEr1UkiA371z5fN3LOucZicdH5Lqe3AUOCQRATsH9qq2cFQZbiZ7LTrB9/
cht6d862lHQQoTbn3ZsewHXqeeZQ5i7hjzw1IgEc5JoFZFh1Wm0mJLMMmYrqZfZe
vsYw4LV13tbvWXAcALNhulnPrWmq9xGtscpOL6qfGitoUZ8LoLFykQ+HkWY/yxZm
rTyVCndXbuzdZKAi+M8tfCKS1CDgX83kNANLns2jPsWutUQ5bB42pRiC5Ng4Oiz4
td7DRvpIMYzLId8VEudIewBVworiH4QdNyfUZWtCq7CP/jzbdgbW+uq8ApNFPjQW
qP5wJuqokUhJh6EkafLULh/4HLL9ozCPR3aEGl8BchH+XlpyV9+R9EdShWcXSSw4
Ltwn+uiqOurIljor5ywcfV6QC14BRwXNzxsYzx2Bx3qK5emgb/nY6jtDnN01Qktj
bpUlHbGTW8yLQoK8LPw79m0JT3NC04II4f322Y3ECOSDWIXWbq9AMRH2IwnNO2gq
Ed1YhS4h5XeVvqDtwDOssY7JazTgoMXQ5yOxvw7ugGFhJNuj7ls6w55AO13U+rMK
RFVYaZL3NdQKIp9EJJAdpRwpWQuKRsZOziuQ4Nc5QL5q3p+dkpu6uydKTTEqhqqs
WOQg34hzBCx6pz04mWFnLP6BlyZkWx5PiwjKJ3hryJyzOBEHU/L7Man8CKnIOhzL
ZKFabV44lMjL2UK0opsqFI1KMFXxh62XM5ZmoSQ1Ry5I7mVQOWF0D12hYQvhnQql
i9S2SWrQSG+RTP+ciqZb7/YJcanbumwzzz9in03Ex4MqwxHU0WC8U9mGgnOTP6fI
1xIUcTEueFyFXR4unRHkNyWaJ/1J49SBeXi8V8z/DFMVxWVKBSAlmtwUOJMdwDI7
ZFKsY9GJG8B9t6nDBiY1UwSqqKG9M0ycr7MT0bP4FWVm745ebOCHdn/RbPO2o3Ao
Qu1L+CQjTM/HEcrWKg8WX4f6FkAdB+TLH5/18DoOiXI2dbiY0lMAHZniAB8UVQKJ
hVOrc3C1wiQ0qNuq6OIEncNn0d7zSkCI7+uN+fooWsJ4IdkeP/0UoqB0LXaLps4u
dD69o8Q2Ycfe8eVB57+Ifa1X3DD78fflFUXq2aWb3T7HrKIM/2m7oAXi+hAp6hGH
4MreDo5UYz/gqUfB0y4NZ4vAflmcIblSPd24kGRba2rGNOcpb2HqSa6erdUEEYzr
O5J05m3wiuZ/L2766vClfwTdBw1UAT5CwHTad9sD0SjJgKSMmgM8J6QNDIeNpovL
Doh6nFwPj6LkPRmLRBR0XM3OR31t0A92MbjNAxLUnK0qk4cvXzkVvv9CejG0EXYK
dAyBAGIgPuqVu0TQGDT+KsYKar//ps3OzRS4EhpTM+UrXaqUXksfnQKeNrGwaM2A
m84pDAWeN5czzCa5E6Zp04DuZha7CwyYD408tFvmPrqLv1igi02pmUICaZAWlgr1
BLNOqgs4Sn/vFJLsr9sdGpDgk50vGVDEZ1AipqlkMbYpy0ZbYXmDS180r9uLRfNx
6WAWXqp9pnSMvxirmHaNWEZ6Aev8VV1xBR/4e63zgUmnOAGTBubqUQxdnqq8b8BB
uPoKcoUvzYblsDIKhQNSMSviPFsDGuN5mtEgBULZrrTYHyw15WY6cQ/kIRQrU07n
H9ij5p3sQNnBiTq9OJSXvJ7w/lCWWBR8Hi2C+n9wj139dCbYGUogR1DihrE3gFSF
jFWreoSVcvKmcfKs8CNKBou7YMakzvo3Ub0cYn/ABe+oajAWmidg90LyQV/M5LSZ
y6HRAdgIpqr4A1q9GEezt5aP64kVPosKodgHbfMe9nuSBzniKvKvRpxOO2unq+kw
5zdDYLLUJa9FGwXl6q/EekFTuC2vHEfvb9h9fVpO9pdD2dB+nlWe+wTy88aWuSUS
dYfRU9tJyOeCyvdhTdGwBMlFO9ZcZ6gmFMars8BXbuBVhFL30xfobS9q/lin6MaN
dzu7sZC9/P5PUzKOcE5rY93NHhLyrHiq0UI6fHJQSdqzNDaK9g1hVkXe+QiRkgZU
TgCeoMT6gTWP/WUuUnZ7tP6nAkg8QSQsAFuUnjEThy6nVrACq28LuecVaw6AzcqW
svDK5lFASBG9ZPfK3BkqzoE6JGJ5OPoKDlkYRGl3btmzciPtqrjz8jGfd4pwWpMb
81ttpfnxWzdsBwkHX4crsKGnuiBFFE/uUIonOooU5AxtTFWCRty5MDXhhk+fI+dm
abT/WQynyY6tKXmsi0prbVMVO91k8vGPor5NvXvFlwAMoGZJHNWND42ZhAxakUga
rkKulo7PHX21hn2uSZaGAb9Ixey7H1s22PbqqvCyV/ypIWyCuUjMrGAmwFAhXS47
s2ygL42q8L8l+TPeFZuVJyAQqT0Q4LV5M7enRKLjLvWxMtqqL83mvDRUlXFfiBE5
v15+fm1BIzIVZMZju/f/n3YbGBmPDpk7co43qH7+2+D7ukqqn5o60lV4899etA0J
5egP3ehGmXdsRZGsy388iXoazO9bfinUnS4/JZIZL1hKlUFO6I0SC6Fjz0FwZvpR
PDrX76SjxWTqMngE94g5hi6bTE5KNkdfyyV+61UzDAgu5M9jQmKsN92aYOQxuaG7
vfDh+O8lb8UAbZkGstwbk+072Xf2Gt0v3+97A1oe/ADyPAN1IrMgc9qnJorKWyR4
U5l0SVSH6551Rvd2DZHEYLYK9OdJmRLN1cPa+aynfzpng/2B+Yk9tRluKJwrzA/u
U87NjaAIR6RNj/DWwlh+tSGkLUmZ1KzkgYI8anxgOC2rFKQzNkAxKfrbOYai/Z71
XgxZYtc+bB/cuPPbqkiuYMvSImdxxyVo/ZGCBM1tPodRokmB2rzfdL4SFK9WLW06
WTe1giKUSeBcmPxM59UJxr0TtAJkZ0SFsaumuLZqcFc5iWygKBGAHVGoQzoV05Om
HptmnNOWSGnfNI0h+cnx5B3Afh9c9LThji+XFIdvjdBEPI3Xjq1H26JcEtL4VELs
jHI2qQXDx3L5RGGkMCXKP4tAJRilDXm+NXoRtBnX24YEQyMX+hc0iUL2M7fppFBT
PzzXmt1tnEd6GG+zpEDnumGeT2T5HarXjF4Cf/J5tqZMGqY0h0wAw9lojIspaEcG
wCuOExOtePsX02ki8LOeNjaoXI5tLpCwEiT9KKrlqD3qSX24sQcywxbAu5MiGg8m
hYXcVsxEFapk3qErjpbTshmxu9VgwGUcLNCpOTWKwh2lH+I1z9URnVXq0AOFBjOV
vNlo24POTorTW6nsebGSl7uOfqmDwfc8rydS4S+qeMgLoarGjo2lVor6JzMztq0X
KIfuMLm/0X0xchymM3btXeLbbab52J12ic8O1pTwTL3Ah+M3G+zJeppWP9/4IH3n
s+F9ABdmlo9OQm2FJN+7h0dFyHR6UcjEOclbijfH0N4NcCXoz1dgBAQpqynhKhVi
WanbQob/2mpZQDlm39MBC8r4+W2Afkqi/6yl8QALNWsKdljBpWSAYDEYqlkbgnrc
pCB6+IdfT27wNhuSGxCl3se7bbxzfXc1EhskTjLv31wdBJVCVOO2KAftkBT3KSPl
Ev363UP5sMaULt9EbGpZyLvNImAL+KVau+4DF2qGOSbL973GTQ1dzYK34QZTtm1b
Tuo+SCm5Rkz4bd3OIiXRaHbG7B1Q3gtHRUWBD8aFH+P/I6yy1CNIIS+tlrX6fCDo
5KnNXqBejMw6iXZBqKlnBYs9/tGspjd3n7ehkP9Bw9mvwPaIBDGgb8rC7XbMe9aC
cfzTgvlyDO4p7Fq28AujjbReqhjhMWP2/VD4R4RUnp3nsz14n8glMLOHLeKpoBw+
ZSLXzPeU3tEBmqIwLPi1/7qsYIxGBtSvfc6YUEiWurd1MwkyeZIVxSKr+pkg6zna
KfmwHY0aK4dL+7w11pb6Nlpy97eCMo8xGd7j4vMF4N4PvxnXBLUZhYtynqb3hpb0
yp4/yBH3dQlQndoi6SPHMHJ+YfZV7IIvhTm6tpEtOpMty4hwpkv7/ryg1+Q6Y7Kl
XtVc+j5Nm6ClqZTLyfohOG6XrGssGF/BAW6S9rfLozITsTrt97JwfbIBvYAfUaKl
VxLPEGZsuLn76I5MOZfpf2cuUKCx2eegyqceH0WMHO8fSUij7CAw5GuwMUFDy5Vs
qqBxDTselIfAsYs4tsMV4ezlJbNpHhy0ozSgVbdkL/icX+ySoaVHZOIY0HGvxaNd
h5MxQoLS95QQjtnqhrbgi6VVeoK62/lU9SYPauiviIiKCnJkPHzbHCTa+xRdyN2x
IG7+R9VPjWGDGl21iHmv3Rp6/d5ymeG/CXU3hKPKbCj+nbgT0vOWpAmH0S6ICQGA
eLNSKn2fcXiqyhDFULHeN5AIF9PHxO6RSVeBmRwK8IZ9voRHyvs533Jdzvb4BtBx
Uo0cHhT/dFzfUIgtV3sPcWV7gBBsM1aKeWKW2L1Ll8iXepkrxb+hdU8eTAWVzUFB
RKZycRWrDsSOjwil9T5NsZleL8Tl1Tal0Oy7WZt0lGPx265ZoMeB9v+pqqwk+/KB
K3XxELBkWLIUCwn8PthrdFaXrhlomtxEOdAaLBDj/3nizrm5qStF/oo5aTvDjN18
bYfHJvSFqPVmUkKwHlJ0maJFdfMGo/tlZSlpXhp0tDpvpWR0Rdk8sx8ZbWfK3RJv
Y+mqTnEiCMIW/P0OzbP6tK/bXyJEnWn5zNNttNSJ+irtRLrbxfah4WgPUpXOCzIY
l0hgGF19g3rc6d1gNfkVMaB1AW/2P2vjVtvNbrtWAsPjCs0iBh6UqlDtsQPpkSsd
MeouePjJ3u66kwe7Ng7A/XcjZwyTNuBfbNOefUoC8mlKSoqyt/PyQhrxYmysKSbs
t5uY0LwTVRcHS1f9a5So4v/Ddah4OB+9p0cJz7GlRKE3ecFseXl+PSidxhRZw01u
kcNVenjdwvl5Ubkhn5x5WUHUTgheoX161mwLjLLCRkbZmmLHL82rnuPwHm+X/rtA
AzuLuSBNpwZGFU1E1K0ksbzVEQnB/UAaKc51cSS5CzFOFm1ZTATcVrfCWLircDLf
7REkSbJ4d2K6o4tYSTbuIJMgaNPOAUcRAcaxU3e2uoHAUeujDwBXnlqFMHmDMzwA
AeblFWfFtCH6VNN/jExZLh5iNtK2ayEW8pvuzplnUb1T2tDTybL/BRwxw7iGqeO3
+uL8Uz1CYNzoiFik7a2atmBtcSS0ZgyKWfGdE9Ce0BeYcf2Es+OPJc79JXxPe8X3
uSBsnQzS2M+FuN3GMrryjy9k2sJkPXVVQgFMMLIafg2rjUP8tUaFmL0CYvDtmeb/
/MjWMkDbUBYlWny9xaxq0jIrv53KZBGRoeUScBOzD+Dryzlqy0UzFH5mZruG5zqp
Xv+lnJPGXwbjA4+9IXsJbc+fMdVj5dSHfv+0YcHfPOHJ9ECVy8WWe8dQ/8bxGOtr
qNAbSNZHc7wze3B9ki1BdUQKOQM9+WayVXZ4Ff3vDCadKTyZnb87ORLsCsYE0gbf
iyulaqH/9JGNNCItCzdB/LnAcwDt6yBKxSdyiNgKAkaGi3pOXf37X/30uKEpoMwd
XwjhwYn/PaA8W6klT4SzHXAAB81do+xAVk3LlJEc1fthJW4F65ouLUhwd1uKZ3ZG
Mo5xqIF3YCK5j44atmvaVoVI0Mj0xr5Onplg5pKZzuqFboCLlIhdvUBDs+JBZkDZ
e/ko9Tg29sEJxtf0bxpu6FivLtfKdAXuSXus/71ItgzwQJE6mai/9Rg8Zwh55FGB
p5ExgHUXyAfe7NVTntGI6Xj5e3DD0sjUYTe4O7SpOugiWuUaBwpGm1YvJR8+q8wA
VfEMdtAk6OWkl4ii0Q/4Wo4LboYHlK6AFZ+7pFPezSx6LxRsdI1pC+NlQYuc4X3o
4dtlsscCjGXlMQeltNz0UflKyM3llyitYgsuMH02pVnoiW6yxY8tSoz2OlAJBtNJ
/5gUs82HUTLnEm/Fjy0S9SMBhYWBGFIidjn53Eh7nc4WXVWT81ILpSpTOWU5H0a1
xBMs4vCaIC4/UIuDbCO8u7A3kUUQSLXvF9VqjtDIDn0DGctktFqopy0c7VLx4rZP
MgyZ+Y36hdRshgU4TBi1hitOgi5kBj2OKRE7ll2Vl7NLPPC1Ut+kByzBeIzJcRhN
3BU/ARrTujFOD4PQXiyCB4bPrJaSLjjuORrSS7gGImAbydHjPMNreYOYj+4VC5NJ
C9arFu2q9yYIc45G2/+mE+BY/wEOxAaiuIWyhf0GYINE0blDSBiZ46Onj0/zmKYj
qU3fRCntWfJr8MG/6KsBsA/UinBFX0xldc3UQ1n049ieO4QXizzlFTEVkM7usrnt
TyR/cltQwZWHa2oB6RHaRy91xS5m5Wvk5oBeUYf29mq6DE67Hh2eeWbKZ8903GOC
S3ZaM19zNNXydsZu3+ubGWSOJKvcgi5OssXPxvpnWY1WNaJwHaBkJyENx8su7tk+
WHLUrMU/qYuBlgxeo+g3XhNrB6YPE5ECRZcePQK4Wd0y3l/ObwY6rZbCjAbLMug4
E3qkZdaxhlNXUu1R1XCqnVDHUxrTlU+eEoRD0mWfH+AB9P9RBFu0DpBg0ZIJ3ph6
a/KQCaw6J5Zarmu/zY/XYM/ziAqQFtR9VpElM8xdIzbT0CdnP3C0Re3q2IMARXIY
GvXFvD+XS5lyHMwh3M+FpfsW1/L1vYVb0FdLf8C76u1fl78+ba5zZ+SmPzCSatce
Wq3yvUVhD7d9tuQOQL3R/PQ7lvsjQseIkEJnU5QnK1Vvp+DD4RMYhBRtB8hwNRNJ
v/NFOw/NWjHwTWhjWetcmrybmvY7RJYO7VabBw7iAfZKCWLozKasAn4Q0JHwlAqi
BqHbcEDjiWMeMjlJY7T1wCAc7eZ7Zff4gOdkf4QRaDC2dz/2ed955KUAzRzDZeUt
TLdLadBpMVjNxMvjSQUhpFDFQREi+Sfj6FaJoLMebB4WtoNLYP1RswWfy9Mbc8Ws
WroVedEJVg4iJ/BVSZ8hU6ET6DXOPmRQll28W+41vGo+6xcDn/OUnlrGIWqnOkY5
6dDT2c+dUwilsPAQYC1tWGCabyCMtUa6U6JS+BzqTAYoh3dKRkP2SfJ58PHPSfkT
kwsazZgsEVhu5R4cIUX8YOoBiKxsXqyuV1WZFUvSuEo3RRoXfZoj+jF3e89AmWi9
dx9QJTCbl4vCWeTo0yBocQ5uMKVN7AFZ+AWln0uvBQpOGjyQ71WofcclJ7VKJGEN
WpaBQ+rzJMWJMI35Sze899JwXi8lAWb+xxt/nmO/583y2QF7LpZ5hvrKJ5oG+WhN
ShbY/es8jjD9g+f2xTzVRFPMsYAUVH2zpzejHiPGgmAWuPaBngK74YlCSIR0RWUy
0iQ1jigt+Tb7Qu213wwLt4ejMvvi4YngOwKF6ayzyD4huTCgmQ1oanMzxpDKu9nC
z4OXfawytG0lT5OphZx6cYsSfcENoO/UMXmah3+d1DqBb4qu6ITqUcIwBzjE1lyV
1X3AxGzR6tFpSEWDmW7mxY2ATr/4+jSeBbXoq+aIQ3Tqw9L++vAIC1IWQTkARPsK
61mEWCaJuZycg/DRmrw34lcFmp5wy1x6F6d0SWKU4O5/IeD0OpJjddCk959JP6Xi
eUOt1Ij9AzenZR04HvakH5NEZfjqsF6LUSKWZT/fJepodvb8gnJ95NL5i7H2IuZc
GFzWHjzCqYzk6hplBi3jpfokpa895+IcnhuAGqvVprH8SOuPGOsEOyKt95LLIJcb
t5WcHrMXMvLpyx65QAFGDBmg8ApaR5em0nlpn4C8cL2MNDeSTNCzzIWXsJlkiC4a
jqSLiWJOYpUpBm64nl3z/OXN6/gMwU0FZxAHrNqiLl2gRU1mYoMcSFAqptahchSU
ohz8aOWiDKhCY7DzB3JoN2+5uRXSyfbNBiE/OSj2by+FP6VMNG9chPXxoGI0NujI
KBvtStw48yNo4+VsQjoASLzvor3ItIp2BxOBPwT/HJkk2wDmHS8+JpxH130pWnTR
b4PWvtTDz94BdDjnj+umgpSdM50CIlXXgNrOMine/BsGlYtTMS1mqPaasC41DVqL
6smDJNILOrZCSWpCjbB6gx+EYWrJ4ijMxr2ciw9fQS++L60Y+9XXSutdm1nX0om3
H9nwCH266Yves1L/bnhM4eGKoIBbHrKjh1Eb0K3+vtqVfSx6Mf7Kk5L7LCPgQH/g
B1OnW0PFCmC0/t+M22b8zo+UG1FXa7JJjsoI61/AHsuAFppz0eCAX6xpyl8Y4usU
vdzp276VkETnx6G47CYHDhXgrVJco5Jf8yWgCHpYKkmpdl6kLI/1MZGjh+RGLd0u
3kNq1wj5t/S3pRa34kN9UMgN6ui5mpo1NZxGpqOt97gh353iuYiG1tZf8lqUGRcX
eUbQNE6hlx+eXJkbjyv0falw6FtA+t+Ub6RpGABXQlW1CFb0p5yVkpwzDC7gGYRf
oGZyofw+0q/JuEQt3+DI5h7V+mXZvmH+Hk0kH4wl3/J234J7MPP0pKgxf9GoKzVY
z6XeeqobgRIKEoMidIO0+9Qh7NUDUs2ahnzWlqs/2tw5mTkU3r4rRmnMrUn8s40a
nhkEM64/xoC2Bb0m8g8gNSuIoKiZG2vNz9DFR6U1STtBnhEv9hazIY3KRafvDqgS
B5K047vTaQ+p0+1Y/dDZXRq/UkPrhJWqboonkD5mikr2xeCVJtUVQDUPBf4O2fz5
siGyZ4RqTI/SqxMeKM4rEIZYIKn6IGjIs/hWJF9UVQZsIfH3oQneA3WMSOgoIqYe
wtOz0+UwiR/bSWng52vrcATMXZGnydNnSGArX2fysIyTnVrLBf0t9ESezrHDHdRb
rmBWLoljdfTIvyKriLtybW5ZFI69saRGBXxWJz+q2FC1hibZBnszatQo/2JakaSG
MggjQSmB6EoVjR6pB/rnGhJVEytAy4anCWIbifFp/aVbGCAeu+IXggyk2vnJgGH2
HHEYeNeV4+BcsGVCVwZBnJO7VipiOoxnf+QBs0jNutWmK69J7FXM23AokoqeRptC
CtHIvX/jaLLc4HoNQ/dk3y9KD+nduKZUwJAyQsuxgoxCk5xY1sBw2aUD+e023HyJ
NMhLBs8ZSSIIBP8M9Xo34oBFKYkPMFgSwf1TXqTw2SXTzCsWBhdAYoRJHog16ez5
H5f/LgVZwdYVZJjI4ByYCmB/PaJz6sO48eFJcdjXN4uqYDad/QB2YgMoqxSrKpPx
3rtyZBiDi84hanX84B9+kwgn/ik5dwif4BiO/7KcpytM7NP5t4OQoigc9SOC8mQO
0QHu8RPSOlz4gakhBHWJffjmMav71aNaayIjWgY45BMCR6ML29KH495XgaTvrJwL
M1MRpKznnc/w7WpOB72QZuLWbhI0fA7fsS+968aVjS7zWtIzM8XndNnb4Ci6KIxF
K+xMREXErNVzjfsr1ktXldOnY/Y6uAG5EoS7dr7Hu65u897bIetyWDgizlDo5ByL
Rcz61aZIJwEAs3qFG20vta87g8klodimH7cocymJjIHeFUx54NmaDAawLwZ99SIY
iRkz234s3RJdNRcl8FjEd2rT4TnZOkoz3CHp+5M0hldxdaWT8EEf9oPo4o95TxLV
KTYKGs+9KIfN9q7HOFPFOp3r6wEhlwp8iZdxuxYcCprW9GKXlX5Km8pXjPFigb4+
BcgFBWR5EacxF3kbD1fJ0eFR9ig+0kH1NIbJpEFhDBNw49dQLl8c4MJ6Xw5ggNQi
70rXCmLgg9f7vRlzZJn3uX9zhk2k+3HvgctAy8GNF1QE5SddSCDQwiV8bXY47vPb
QNOibECAD791yGL40HOe1FGzF34NRCoY/AB7Zcih05swHfRvzceHPrCq+7DjEXY7
ueAUPj+kW+EFfQc+UEyjdfhpqAPFTsKB1T0GIjxrqhxChG6dKQ67jPioUX0InMxH
m8BQU+jfCe9twYOrtVVyMSZCV36PrqraBajFfV7sfU6QDSHrpgqDD0kY1EPFRcSY
/hiXS5yHta9p4fxueIW8lqhtgx3RzFqrGxDY/L0JLLSCRjrJes0cxbIv6JXPzv/D
M619GqGa8OOMp5Ma0F6AGBxO9qXNQy4m9tus1JVB3GDxQ/juYZeirpbbq+2+aPQd
eel59q/pF+4/ZMto6aeFKdSZ0NNUcsD0CFsuuPfIO0GtlsS0g+gA1VTc2hrADYHO
EvFFdNxDPM+zYMN+RB52SscCj453yYurIhcjdGXgErhrZ8D1i3fXY+8y26DBQmju
TBEaKpFSN1o9Mqo24vMxzUNay369YLTGaE0UZI53xX2vbfm5QMsZrxFjHLeJH3ev
tefej0wE3MYr8cDwVIkFUSMmcsh73UTByFgKjV4IX36nMCO5NLgyA9aNdl1H2R27
iCecMV7+xTv/WAdB47gyqJhCcuvaEku2rajVR7SlOMfSruGwnsApIpgd/2mxxQBN
BLBE76EMzQzglj2UYsqDtH6wWoz2DHZ6u2V6YRJfDZdQxMKsx58pAYBbIez0gngX
DquE/yywDGMEDarsBKnrCbsogCyzMOophHdZwCEEeJNP9smKMZJy4XLppPm7wMRN
ST6Ax7EbgaF00GK4lj24n8jDwSFwUhT4i1Nyoj84ZklVAXq04+FHHx3W7+6dfOc+
q8nUD5WOqLuxfDjAWBnuxbZpgM0W8VehS13UMtK71iaaaK9yHEXCfz+DYz7l/O9j
z2Df25paMJeVVUgCK8eCvIanJO9OcVPBM2n339GlGt/ziHPzMMMgc4GMvq0x/Uwr
bl88LKxNwcyRXiGdF7CuYj4ymwbYvJEXcpJ9V1EGYRB5TsbuWRdZPGaXoRBStDBM
4I9SOnbnrJnvYvaYqeTYP7iaWr5k3sVGqyO1ID80nmE8tTihb4F1xuDKSgA5OHA6
OpQO8Mf/mQnlmNkQhrgUGjHPCGXEGWObv9UYc8vr9B/HfNLAbyDqkcDvM4XKXQyQ
Qg3SExY2QQyU+ojw9aO1xA6/LLqpviUgs71dTCcCDfnYNqyAwfRdamEm8Vf2opED
AHtMaEmWaOpXsL3xbGh9Wn6PhDdYZLi52FlKUC4zk+1S+KA3yZgOxf3to9/ZCMtp
d3sfpzTpRwN5/yhP/eLA2Ms4iLtovkL6igmi4Xh+2DMDLv7dTqYgL9MoUnxbv2Ym
pValUXope7Ma6n477X023ymEX+M16cba6jGTspuu20ZpHcCDNl7095w3BZXNRniQ
3MbmcVYLroOZROiiAaorviCAFKJhclfkD2u6qDOG5AqTFkygU+PZemO3YPW/gd77
LqJg3e5DYj36Z2j66fIRt3qpZFmX6ZID1TuynQPku7UIAk86SJZgyt9KKiTbJXEC
+2pmsXbJcBAQ1h+s53DFRfkpR3HG+aKxzc3Yucc676pt770GpmROAeNUHaPs+EGo
VCFINsJW25vttqAQuYxjkGkEY8SfCaEQmlEh6+GO33UAcJWElM8MZ2kc9qfjFjje
Mr5AjOHXGwxFLxjdKM2dc8zGDL09OExuHpzBFGdhmNhwGu07Z7iFb8hdYlln3MPZ
gybmofMmUe1yQALPT8KDu5sgEMRNBYX8hB8MT2qxVGA0keSCyZRJAAnk55KbTfio
t3mVzuCBXq8v0246LctiB1CWsoDuK2HPRwTlvP1AGczZLBndSKzP4cIhByqYMqK0
QZAeQpOqJ1SWcNTNY9R/+T96sUWBGcZfrKK+j0IW2FnxQmcSvtDw0P+FWSFdBEc7
QSc+s1/2Yqrt3jupBaCLAcjqVbHNgrIWD8/UrDZEIjqhR0dfuddAWms9HnRhRrpM
c1Lrmd/CSyEmYPRMpMdpD7QMb+A4kBeo2XnEbnOxYYE4Si1BjUJQh+Vs6eabUhLq
5hOf7rCLWdvvZmlP7yADSN3OLTWEQFR/6ypiFNt81yq48AApV/g9io4pZ619pTd5
Zuehe/3acPhUk1LDc2KzdSQt/JlAgwaJfTgtNy/yZ1F9IPOsovM7DEFzSsmxcfiw
M7CVl7+Uj2ymMoqh10vscP9i7Iep1zab6vDpzFoB0k5T8+6yGKnxLvY+m3MA2+zv
E0OcWZso1xU5/j+QLOa63dRMIQuSyfEAr5nWbmMKehjPt+xYueL2rhK9PviKcu9p
isBfWYg+Yezwlo4VSo9RJWusf7OVDo4BfTayfUNFEcrFY97YwsX4extIDKxmKw7r
MHMZSO5adYLldXiN+uJj0ePEwt3g0s1aj4588DPCAxMPEsoxeU6nOubvlZurYsXl
r9YcJGa4MUypj/7AUm5prerFzxl5gzS450dT6h9q+TpRKFu5U+HzM9ek4OutJ2Ks
/1r92sJg9IfYVetCnFU0psOKNb6H4KA/iVCjouFtHdkAlNe97YWtsU5UtBYn76k0
V6hQg3bXzbJsYXzXsJS77jxxGE0V2J/1mvY+3tOByTPD6Atv57J+k8XiLriM5wuL
lxVShAg921a9aUZpCLiy3grBZDQ8Bs6Tmv9nm3Y0dkFHIexMN2Cbgs8jDx7PCxWK
Rg8yd6PDzE1312lYPaaKGYM+0pl9Z7AFrl+WTsU4Gzv25bI/v8uhAHWYsWs/4CFP
ZnO0hbwdLmOtsB1AfmK0hKFNe8eQ5e1kKq8ll8y9666dvdbm0RTPb+pHfahb4bKF
fL4dKgUwfrFQCRLXeYqr9GzyfAfcQ9BJrBrkzz7aI9la9dd6Jm8OYNPLvOzWuX2+
hDkB0+PtpxSaoo6cpW6qkj8IILmdsQxkS4oI6Cdz3gqVWlGz5Qmkkca16rg/l7Pa
summDbrQC0Cix6HH57BEsGLQc8LGJMDIPfHJfehr5pMqyboJo9bNh4xDATiIiwEW
KVY7G4PmEu1aimMAhFayTiBJgmIG5ZdonnGGt4qwUr8IUryUNYCUnka07XNjSzl0
uTT46wd9j/lZm3w/QQHM2q5SySh6zpkYzb17duTnvrmd5SSR7uMAmiyRiNqXaNWZ
AYHmsWo/22Re9BSaFTjVq8quUC8kdRGs28obk0oStU8Kec9uKQxpMtlZZG0Zs9lI
lvv9ohLsopgB0ovn2ty5777bf0BOZcEQjyeqKN3ceC9fHat1sGH7KmjdBL49sBi1
t/S9nH769bEcFrtlIXLyUdJ6Pj6tG23e99DdFZCNZ90z9JBM5tMGzWpQZq28MdCK
7WgLgWdFtcVZqGNJApufflkPwk0TxEbRzj/yIKkHtrfXA2RmRPLd9a07ZcFilnPD
bl9iwvW/KphYzFv2Z7EuxVM0uNxrp82DTlmzb7NlQyjqHJrbI6lfV9H03ybbs1qh
ZZxsER4kXezyjOufBjujuOpGcH4H/kFX69RRNEvDJ29wl1A4bPV771IvnbVCWJLq
m3gPbrpW+ooHMVqe9lDU+OMDkbR+YLg+PDYUilXO3ci20PnOgpNx62nAku+45OY+
OkvwXzO7TXRVCtbCRBSWhtmNQFQVQI94e94kjoqlpcyLlC82cnKGOsU6w+KaLDYY
Q1MChksoVSZQaYeaYMLMQupW4U5rk2o606kV1eMmnxXbXVk5V8sgsdVPMXHFl49W
Hu6usa/W/wSWkHpUi2LVHU+cL1L+IzLy7DB97uDa79gFX+iQ4dMwryEEYvxweaES
9+X5nJC+SR1BP3wuher65Af10PBeaUdox4Whno5xg6fecnws49XrujORkogLNRe6
ROm6mGd0bRzU2xBg8xY4aWppE91UnvWWy2hSwepsNeP8zVCDPQUGQb8zDsTxB/A/
9l6PRdUCm3xtUTodiGCNPvmI4AE9HtMmdHEcp/POiOm0XIsunD9C282KnmAn7vwx
9lSlP8j79B/40DrT11N9b+/qmu0HZlvcQQ6Vpin7ckDIBTqalu7FUOEBjib/SjwA
nVpnpCBz7W38vIeCne6XPsXEa1kBfMGBNj1LCIUye82rwyewCIssd1KE16jwCEXs
3cO4lJ7Ed5WvGVkMUl+Vz+QsdkY+wkMn6SJBNoIxFdqq8Wuz+2qjhc6dW7p7PcDz
jDNLXCc5530OM6MbNnPWBlqVQ2LQgY9nboVmzBtBwCUekMtBZGW91BbWQDAjQtmN
Jvw5o3Fc5Sl3x80elkaL3dd3be1KZ0xbCzd8enJEn7qTGI4/GBO1SfcMKELOW5Wl
LY8SuiVSzCfHSpsA6JlWXna+iuvPgMXBPNqxGpff9704pDsyF7O6yZtDCdRR2nNk
S6d6UoRJrQOkktOAnn0+W1wdVbrKJODMk16kZClsorgghYOvhemH5aA46WcUYgYo
q9eUc5yi/MmnrRb8zX8mVJry/3o+Q/nZRdRYmC9fG0dle77WKlbRg2MrGqgBg1I5
FNoOrozVQkcIcsWut/nkP+97LgLkp7JDTAHrOE0+63nseVII8jIjiuYGFIkdLmoy
w0K3V3FCYJcl4hs6Les2JN7Jp7t5NQBffxXDRvbjQ6SvWH9tMr4wvnahx3Ctlvfq
WhcpHNVq7sD7tJ9uX5jwyYeWFtGokUAQRefbas1hyOPqC5qdnxeNmYTo76VNUMvn
o7tUqQLkPb9M18EO7VETsr3B1dFz22vCyOWUMUjRpOynv7IGaiZ//Q3EiiJLqWoB
90kYLyWjAuHE4EczD8Q6RHgzrAXSpOTozqPVKhOCTu6Ut8Ei6t2Got8E9mbOQ6a4
DbaEuJFuToLeDBY6D4Qq31dtMHx3y+y43ILC0vdTqPqYLzfQiv5N0PM68KG5fVfe
xjIDeQqN9qMF6GG2qaatxtb7yVSfqVYvHD6mAzUiUurGAXPTJUxEfwxnampVbv38
8MUQ6bTRrS+5O59RZ46g8GtIeP27yKmhT2CgLLsHwTlJvx0vtH3iG5nD1bC2MVF5
LXvN1gURR+99D8eWMlesjnuF9YO/ZrGE56S9HTH5WzefeJXp/yuCM2HvH8wTxoOv
fXt5UjJJPbYfhyx9zsL+bMw5HccDmNHN8iIR97QQQMv60/RUCXc/r3yOF3qnWcHD
nN6g0KREiksDo9aIlT9MqWDbaJB/bsbt0mz60Uv0+97H27ne7mkpvhHyJ75QjtQl
h72cWTJEDzj0v6mw99Db6X7BArS01AccX10iRGZzCeKhSpHopvnATQs+YbF2oUrZ
aTRPeYCpFmXC0YG66k+DaHZ4EfklycFf34NOrjnJCBVuWK1fC/2m61oBHuQ1bXSE
7cisTdvqyOe79BlsrHpa0c1sm0gZVz9FZGan/TIpHgVbOJh+8Rckw+nezHFhxIgo
geE7MV00luHNthJUTT05bbZtPv4K/Ak6IhYdljuCc2hGPk5N8OpCKGDdWoDPAMXj
OGUsaNPTSqQThW9uB7ly+poWI8uA34/e/tvFPu6Xtfio0ihJDRNb7Dob3VnazVai
j6sQXVejA7ruIlj9u826T377PHHzs4Lka0NAvVOvgxFBoa5ixDzhfShRblb18slg
zclLuvJ84Vh8LaGVZb8jluEqGKafemCu76y/hcB55Ae8SToYhbie3xnUUYSRvQI4
JItJXM0X8dlHSr2wAwWPMZCv9yLMwNuZF5hlpOmJ10W4jYHVqKduFK9NDWdTb3Ju
FvqhMfIeAc6+rz6AvRMK/G8RNG0/mybVHPo+ubZ3q7IeagRodnRLKU+7jnkkxE5q
44mE8CTSv1AvSDx+21ygPpWEHUlZTm3kUEY88EVYd+dOYGPKP/y8A/grq2FXwsDY
GYy2lukdb4rWwyqb4QlCJR6xXFZW/AIwhUwbU8xkunjsX58FJ2yrsoN0RqH+5KOU
yn6FFvXg+7HyihjqYsh1U1uq1MuPXgqtSa305Igp0K/nCEagym2tMTruEJoOz2fF
P20wouAgr9SjwwRGwLPprQToarUefOhcbW5NWGhLjGGPdJfG3556bFXWLQOEu6P9
iDVraqetidH0po5s2lB4MSUmKeRTCrZF0MBCv4Z8K8YVSlTZXVYzsf3pXwSinjWk
idGjQvi6qZebwUVHoups5p6FZArOvg94aNf1INYB6Twd8FzlWfIgOpO5eKhAobxh
tZdW63PRocHY3Pb+h4SjoWOFUuRjX3yBQfthdo+2W2bUJa5Qhfsi7MXvpy+bCYuS
9obtW8bNgi6X66jGm37RRbVTZcBx/D6GZ0ZfiRUVvotyVEqGHCtAKuCSIrPnHx5s
6+fCT+VGhegUldQT+7OHEa86WwBonKTvnWuGy9dbEsUfIJNZNlgSJKD1+LWC/Axe
s8qhAlL468KDiv4xX5MdD//yudZD5krmlBdZOh03fKDBrQCIGE+nyl1U0fCtONH5
85uZNLCU3zHGrWzw45sVcgXlXVVYtwuuKhdM1YcA+KudnhAPks3wIbYKXVRt2dQy
jYr6kUGoDPKM7RtmsaDcg1QCmLI7bzauRZsliSaTTJ+wqN8JwxCa/2MEAhkMHJcI
n/6sRqK2cq2/fTZ4kyxQjgC9EEFfcKGdXcX2QCSE4yuPDUPeF+QezisT9fafi5q/
PYHXTgEvpM9Qzrg+8dJaKh0NwveQdZ6RRPqXWq2zAgLibqbrI31f1LE+AJexbla4
aVO1lak/LkKeKxnBZhEMqCxx1dC5xKH15mCgQ+sg7JeUmYNCN6XRZNgBPPyvUIPp
lwik82CQuR4GgjK+iNs0NsA+6fYpPMObAanGuzFW69EU/h7DvM7F3nLKxvJIOd12
kVcr6mAccFPjUTClxkOyTGoRA57aJxiBJift8evCkGZ0BlgBmluUEjeo6HjavaY1
+aqx8V9Kf6+8S5jg9ZI909MSuogYy4STsjpPrrncUAXgvknAFp8gROjPaq1KHThZ
PH41rTUmMib38frAzGNO+zLKMMX9hM6nTIIc1EfrlWC5nfodD3DSj0un9pV0goNF
Ocm+FdhOuxszS6pp5eHOZlQb/8QZpb8TcFPiJaXylSkucECIUUKet4q4Z0+3TZkE
qyK15mH3gsrmnHhDwv+/ixpFHpeHtuMjm5Zjp1M+LFLsemTFicyCSPrjo7UnIdCX
YKg2s7rLmRY4lT0ZSDEh24jFl8q+83K0acC7bxzlKDCvTSQvRs8fiZ0XMiIhYm4i
UTU2qQyjxvM2lXeV6tlgLZmwJBmL8GnLmlAMJNmCiXDRBZRZa+tAS52jFg8Ekjyh
lm5bHIXx13DECpG/3mUIRMDfvt6gDQ/Z0e7+xSgErsboaOENUzS13Y+eOG4PkOKR
1tn+4ggnYvMtNMOAPzVOjP/S+QKm+VI/OYRnmGa7Liuejsg+mjeJCdHAtqZUu3OM
+/0nPx9WP4pvbtOkLTsOZ/cbDb1kOP6QR8yOQjD56X8b3nx8cRe8veqjaWJV6rt7
nZofNZowid+7R4C0YXk4FYkFDN9F6mo5P8nHJPdLcYCIzJpEKaLlr3c/os4Zb839
6K+k6MdltrKbSOdqC+P1cuFgA6BEskf56hsTzn4YXz3VrivV4V3PfWQor5e9S5oG
umyWiKSFid0WAl7DTpHG86n3SyeWTIcVD8q2g/43PrDpDU+pxXK9ZWSo4FMyiBUW
wjrTO/SCrmU/1Do1hn7PaFrR/JErIczgFB0QDAHb1tuCPLafiOXp06tnAgEZe0kO
O1vvNSp4N0FWdvXMcMb1sNHu0jl/NIqS/K8hlvN2Yd35b6L/OjC19tpJ+vfv8a2E
mN+bpCPVE03oeN6GqHHWgKnY2RyM1+cAG3zPCio59wifkQwQblfzLyOnuYqhtVf+
x9Nz/akkJDLS0gNQ16/EW+p57LAeCTz+//RmMIX0DQ5KfC5DrPUeTO/4ddxNpmR3
r0FULAFglkG4PMpfgbNA7xW3g+6Rtqs6cXtX4ZmHHg+zrIdLN+yi69vRYuDhwfrp
ogXQ6usKmkjUOyV9+RGUqzAQWDqdU+t5FeAdNawYEoWdHckSGsUNlrmxzc1Hha8s
dYvwnMCWjaf9PboTaqeRVTk2dnw8brrwwSMvM5oZO8/fD4EUdksadSXfEutxuyBa
/LnTEUUPx7pBfXtUM7Ni6HrJfSQ4YOP7MHDLyD9M82tEjKjGRelZ49qDe4C3Qr3I
zqGCrhXwqitFWT7At2YmsWW3HSXBxF3fwN2ZgMYd+5DBAi+V46SZMEOurNiioQcC
YQNsu6cDoHn8L/XPaud2Al/NdOQN9/5g9Lih2F4WJxhYd4MMQ82MVFU4JP7NxJoo
F8JJYuVCDqA/rZFzzjSVVWANxCrSMv+fjGXpxN4lvlI+wFzk56gjVNieU72H0DxD
Gt288zbqVjxMNUiTtXA83cfEGZu8I7xOSM1FuVlwhuLd/i/e8RLbU72TfuABTm20
gFh4vNxD4zleOeFJr8pzuhciawQS+HmC7OeE6y1G71vcsrVbncBNk9cLOqkdlgyo
Z+u67hAypaccEoFlpQmJZBHT8yXMC5UNkySLNmocKpiurd3qNxLftod4a5loRuiz
M9T2sbcWMdh1uP8uhNi/fk196B2wBOGKdsWwauODF8VH0mvGqptPn6BkEIJ9viUR
3BEyVXF4lGEVx2t6ICf3lcSLLEn6PQl33FzMQEcTDeBZ2xc8rymZl1Ao+24+khhf
QAhk0XWFd4JLpU4wzG/cIKTA/CkqS5NP06R+0VoDtP0g6hR5Fi69s4LqSqtc4ROE
RJ4b4rnUpjoJ4LzcXSmrjdZuGCDYw3PSBnQCQW/KBTHIByP0pWuaMHEnT2JynGir
SnEZyni9roT96cM7jBpqhh8GgGpxg9LRvf7qcZ7L4rTqvjbNUfIeaCO2q+t7k+Mq
OckcIicoCCZpjJudyeNj7kfe0XX19tgdQzFQ9FOLbZ5w8XdoOD7OnfJBIWrI3SCS
IwPEU5hZVUYnpNL0kctXchUG73cuA7HQrmcgfxxZgZ9rlYfCJ5LYgFAxjwl0C5iY
q7S4H3mBEhFP8ZydTxJB3olnsVYIgOnIw81xRuNKF0Rcl62QpHah0UI+OH/ZeqPq
SqnMtNcnjeZosBUCZNgZjFFAzrmBJRZf0R5i+IQTKala4mgLluVi+0YglF9QGUmY
xtOet89iFcBxmqmhjYspjIWKKuLejtTrib583szedfNP0jkfOIXBdgPOulAkS4yL
vOmd8dEf1nBrZp6rewUJ+T7l9zxybe7+27ti3HS5J2P9uQCzhDGZkBorI95UDs2T
9W+EiTPdnYoiJ37Fvu4fFbYWOm4ZDnTrWjczgJjKZ2NosrAQiU5kRKHsNmjoA2lQ
UdVtOzrV8g00XYXH6tspGsnZ/QpnXKq1s9C2Xy4NqzuevyRpO8m5Qx8Wkm9k6oZZ
iBd2+ePAVEmYU8LmHmS/T3WckBwNY0bik+ZdtKtjyAdhiK/Ty8gZLw/bnNMLmZI9
Su1Jb2HWb6FKSZyGIMCOG/6AIr6z65DzGc3Ch4GE22QuGx2nn4iWn3XnK75sTl52
9L/V5oM5uZ3LoTU90qpxsdH/obPpgp2eKMILsChzFCrR6nKO9tbh+gFWk0mxn0N+
ImBY7ypSVtl3QU19veRQn5C31dIt/D4Y819jQ9c8EYL38AMMCKrg30AH5Qu7IuZo
p83NoUNirr1cUFVG+Pm5adcvcOBN/iVmeiH0ORh+wIQUQgVvuSiu3fQUPkRhZeNw
WuGmuOdmk/bTO++jvg1zbjlpOWDaWwgbRMSf3gieDwi9Ycs9R1bIHCA8K0o9WaLA
TBlG4qDrFfkqL4+TGh81Zdsfel4WFFCOZUy0CkXmLyM8H679RcWFcVrpXBHQNjjt
dTn0RM/gfmZneb2mltQxk2ySlPTtaETrOeCJ6vddB9+BqcHljNqz+4QodqJyFsBc
vogT2QgM3P8voew/d0eYlpgnWtUXN1IpvfrvsB2jMTM5if5nGyBCQspPUejBY31/
tyiJuTClDn2gAyTQJgDIWrEEZ5rEW+EbYrHjEfYLjDB7i9jtbpokvwNX0N664SOg
DWcFDvrDCIZhTKs8tapzk0WhHNhkUon4gJ7uEoPk+MPCY0+hqcD4NYLaKaK95Kee
Oa1C6xTZ73eVa2J0J0H5Q+7RqUuUNRjCCrTkulGJ3fIJhVJQI6oqiMMsJ7ZODNq/
qY3TMzkBv1mfNWQYJfwnYoHW9ZHOhJ3MbkA4byw8FTZz5CIH3XF15Gfiwmt8W6qo
wzz0gxEUKYD/705ZwiOPtjPqAYjuYhIUQrO9mHjJu80aJdQny4V7c60ogrYqef9E
+D31DIWvIk8AdsAeWwm9I10UptWfOK31JAY25hFKiSm2zW2Xz+9dzGus+DtdIL+h
MVjmgo3B30suFAwso2/UyijRbCDSM8hCPrdpLAhdzSDsaSKjhBkY9dEkBZG6Axec
BETGbLgFGyPLIt1rHp9/+U6nxTE4RFRmyGtiGQXp6vd5SQezdz7HzK9zDHmfMZUD
+xxWHXheDxsQwqv7iEpfm5WajvolQ1G33MUELcVGgoOKRKYvK6CydYHsqmRlrI+o
nnyOAJINSrgiykU2aLHar1v8+oBKqCT2czOy5rWUoeKwhU3Smgy8Zp8mPQdJ/bos
wwX5Y/4l/QlZYRCepF+XltqZ+C+SBjqzOlZ5mzXUDVVZLnId+A5JSKsln2Rp8OOz
OMO7t1SfNtzDNJ3nDl6+1vb4yxjksKV6iJW0vCYyoZLFLB57L0aDg8dJpapwYqdm
oWPdBdgDOxaRNmORjUsdUwEjI0In79TjhZBLtVwDVAvYr/m92YVz3U0Aut7S4h+R
rFxsoIBZAN87TF/+pEG/XVzcrqkXZQNm3t0FkdPa1MO+SB4MzYcL8NcjpgYSDKDN
r35rnJ0eoqM8mzWqd9h7EGRCh8T/IfuO+06nl7pIK/6Y1IcgSYTkUm2zYXDAk5f1
N+Q0B6nr3gUEUc+PbgKgojnGLdK0SWGuIVhCzIT086WUKassYDUnTvYthQVpntnM
8oIacv5Pda9PaDd+gSVt3jsCOHMMSfgXV4ao4U2URmJs82P4b1fLabyZ2j25f+KI
INCpIusivJtB5K+iti7vLWpNQIRkCPkPhw60QZ1gip737zNf+1HObUKG3Yy4hXeO
m0imsYnJmYNRQOoL7dthpZnp7pivv3GnhU9iJpojfJ8VFqlqTbA7JuJWx/yg7Atw
dtxQw0AfKWwdZ3eXRCSl0LcmwOpShBQteF+nBoNlRBJJ/sAgCK0qcBrBh0yfVuE0
OslkKNSNNPFsSjCy5kYqgbkW2FDYDTD+k4y30v8UyRjcwvSBcAgtjDVilM1i1Vn3
geXTDNe9BD2vu4Gf6edIW4ZrYCy7Q+w3QX2bifn/y3O7mQc0WmOYrkzTx2BymOSr
U1FQ+TdZRDt/pDIkBZkZE3BVaQ/KfM1IA/PiUF7rtOhzI9PfqqfwcxeLfKl7L5PS
Xg5IsI87zwCpUVU3g5XMkVC9na0k2agM3ryON/ukNkc7F8UePVaX3MJrD6NDljw9
6Pncrdk3UyYHJmriZL5icTYh9kuLSpo9oSLDqfD+k5M6dBxdfqURC7CtUOMvd7Hx
oeD/Pt/SISHW77/3q7BQRv196vNqpq+udJS76iUKGKvoPEOe+Ji3Vzd0sCkW/nLv
tdhLvEQ2eum0XWQO6uoVlakHPMgaTgojb3ZBDzf2lSwnT8aZU7lAxoxO2OVn9rqz
TpLDbL9EuuG18nk09s8OwjFbjKxGJScjDfn1ZDWZvoPpMbFhoxw+VHIoNEXJKvLn
YO3WBhMmGQieU99IdYvs2u4xRIdhSMSBby0WT4EP+VOlsQRwFjsd4iJaCafVCrU1
gMTlEh703HUbxiIepcHpsD5VTbnqjkjpN1B6WrghILnWlDvE6ERXK96k4GGfdoJd
rG35lHM3mE64MlH7EWoq5OTYGWZNRshFg5ME45FS/8cyt4Nl9+V3fsPA6ra6D9EU
6Al5GnZPGwMpCZARZ7uRRqDfC6AjqR1zN/rf50eKULioDC3hwjsU+72ciapCXtFv
S7fep5JZUhLd+Qsv55wdIXpNIvFbklhBDRgiMtQKdoSPHPQy4A/qOTJhsiQZpYXO
xDZaetZyS0jLb8IX7hMGYw24qGewlcRosVtKrpyiuasjxyMTL27u4IviCJFz9Xto
1zqNTxrytPrpcoL2nSteOX+Gtz9FkgmVOybiAyQqwxzWiCqEEtrsHSg+iRR7w26H
dmT+jEnSrsU3XtbR6R3j+ZdRyMOIVnnAH7mZD4eKX6DjaQ6xJpIniVjF7v/RTvzL
MNTRa4yL1m5nAHPzogGEA7Gz1ErcM8A/ZFMYk8BLqlcmFCrcol3Y1up66Qyo5XN1
5RACUVLKuDc0XwS+7b1Kp3wvsEjE3k6oiJvIuZgs6HQuWVljkJSXyZu7N+4EvpKv
8joGnQScJvhAJkv9EjbJ9rIxOwvIB5gxRw2FPrD0f/Zo1rwPq/nBeVTYNFTiey91
vji6leickdIpSB48Qn9NleI4JdzHmikhSzG0bdzgmi4ONIC7p24vLmuKJhNUfyRY
hza7+b84jtxXexK1KvPkG0cfnHdQWe3nKECSkv/uQ2PIIVKZrMV/EE0MZaEsbpWb
3MX/7nr3mmI6az+5yBy/78fMMSvDq/G5X1SzzufX3L25MZv+gSkbaDsAqYTogo42
5l8Yx4Ly+UotFEbF1pk0j0z+XSahjyY+Au/PG6vnDPAAJeWNGNTq8ZhTUa6WstaA
nvPTB1+LZHYWkzMopT4spNGwRlN3tiMb1uVl47aVLj0SqA61euL5fxv09QuoJsKx
81ceUCGCYeFXs0zf5bt/vv1eRQPnnX/dh7QMPnEq1XFV8uTHBFaOddFGTWALoaqE
Tvf7zcAHOsvGQzxdAvCE3uMOGYBHbNjIDW4q34rX8Tgh3uI3MVvWBe13ft3Pi6y7
XTMmM+p3FSXcw/v1rVkBSX2j3VqJQ3A/hp6zRWiZd3hMiCPSfDhuSqUloLTmdzGB
LKIMUwkVUpyGgybrkD4RI2OdnGjxi49KDiRKd9+Uo3e8j0snGoNZJ4WWR9lUEfzo
uNvAWrFAyXZMo4ynyhSrqnUDDjEM3pxZFGhThflztYBZGI+oMoXjH5H8We+FU6CR
Gyctcmjj2Tji/hI/th58eFdRc+8/Rj7LqNYwEWNNt6w1eyauTgViuvwsGfIKK3RR
icifbDz4FjK8In32OXinUqCCfIKE+K8ArEzZi6BdDiPX5OYM4l8/J+ILxJigjHUw
69EpvWme7js1t5K7nf0o+tXNKZQtkOLEx6m2bKNIl/xZCH1urSeIgT36fu6ZmBl4
PLrARub9G6U1EDM4UETIBOyFbl85ITrMZKsCt6/YzeVeYRazwyWi65A6qKx+lCu8
eQqjUcUksG/jO8W6387DU7+3EnVbGJ8fIRD8twcWrjsq5a22HG03QfITK4XY04JL
27IvIgmnM086sLOGLrMhVJJHqsKcra7bgFHGG5z8CSbd2NhWELf92DCpuvusvl+Z
W45vunHntFL+H3XZBULFfIqENFuMlo9CjMQiJYm+tqzUYI1/Mw9Q4lXt4Yue8GlY
hI9gsoodmNIF7QFiY8ZnR5SoiZ3NSsFQ09Ciz/KSCMT0IhtUJdN1DuZR+r0WNd8S
CHCadjKLG2wWZok6cNW8HgL4P38bSuHp+aXY/hwyN6aBgs0o04uLU0TNOI0gcWA7
rOmohvrkGd2ojY+Ne3a8UwQ7DCCkWzo2flYbvLvBANI7a2is1VbxMq1MQ7Hv6xr5
3rdAmpZkqN7F0DM1HbchQdrgOkgbSwrVsNdSzwUGmZqq+/m5Y45MQh4MLjbwzKqK
T/9RU1QnI9FJwxVhK3yDCCJByyKmpXKRlnbYL9fL0J2RvpoXElYMZK7MtVxIoz5r
vU9znBW5+/K5RgddBGcTWyBsAkjvrB0gzaH6n+t/pizUkfBp/wLn7P338RWGTLSs
VdVLfcA579pvNSMekA8P98z6YEnW3oVadcfLw9lU3U7rklIVM7SJnv/LhfwzY8fN
PJcNvEtFwfNci/c9Fy5u54ag36cgBcqHdxkf3RvTgOMDGdc+3semzISf1XTf9OCP
bziMBoeQzxfbTmOfeV63xjSD1cjju84KSEKYSOoqQ+qLxgzOH93ezm+U2MUurSMG
n92M4MN0McpWD/KM2XOyHjdalVzJaQNX4cP/qBHebokXpFUS1OgdkoUlr6VjCQv0
PEXwr4hgJV/L7IZLLhpF+AA4bEf0IGvopzARxrMfJ2ruGweYEHT4vEBPKZ1PzgpS
xA42fsiWQVkbqESXVAm7Wvmk1L3qfNVcKmyPbRqs26AlrbW6u1dgZ+2tVwF6NTw7
lnOotdsdgIdlCEk5y+1lLT4lGekT9m9Yd+htF7eZyXgBnLXXwUuBti1ldzwa1W6G
W+qlZMerRzYHbQbMA1Dsug4VvIDvI+DS5AkssU1zf2i5MhU/v0AYhqH+0BExxEHW
QrS+5tb30IX8Sz2WJRlKB4YlU7D9EWzqbC0pWOScruJWAn6Sw1dcPCuLuSiVXDXm
Q7CKNudHVwiTCBSqpGQsBFAfwkokyH+jm4WL88/9yC3jkHbrMQ0xZOO46QEK7oUb
bNLaqk+Orhc9mH2ayH8ov9YdQTfBknomTguy2en4B1Gx3Y/69uZAvCVCGT+w5b9/
WjTjOrZCEhp2zWUPBB5KaO/M0tZvy9bCUKSFTf4LE+X5ZrSCdXiZAHr/8Ez6dx2A
E4ZBUKpED0/T/DqxbAa05m0BLF/qM1JqrhUc6qOlleo6Xx8VxDwrsFOE5OOr2+JM
YDCWQNf2LGZ8YoChb+5695pyjo/PUm0Yt6sk7GgtZ9lGzN1cSJ4RpitQP46jU/CC
xTP/wqdD0KnH6dHlHFd05Dp94d47JQRLYSd+hSH6INwxTbfYaANbmdxMib5JhA3i
ndxS23IXCRp1y7fsBGd/Yi/E8U14+pvazmB0Z8zYMzUbFyOc293OBJ5XloFb/zGn
KZ1KEQHoaONezoxqbJeoqVpRaATEiU1CyQKEQy1EOTGyzcU1WdDgeaF5oQgwgw2X
2Or2Uv9fpUyrCkqEoOUZlpcRXYczDmF25s+EmsJCA2X/B+OyxNEj/+YHkX1kxass
q9f2an3Y5U4JTV4am4D0qD1CUbYtXJ3xCidE0mWwA03WnSXlsLHcQKPoyEBscTVn
Otw4jIMsF/yuusDzjV5MHT9TVydAchOvfQt+QpLuesyhURtXH4bsxGKwpZZkixwe
oaWVIL6TB3vXApM8HWxAxA42NHZCy9sidOnPc3gKN6UeD8ft0MSAohDNZZXUka8j
KiIPUknvHTyTLkZm5vJkqa+1sC4NiEgmxqNtwiZivhaQwsSkrVDIbq3OCGiK37gS
jw7lceEaW85NgyTqKanUDP4wvbcC/WyZ1NTw8jK6LcTl1w512xz2j2rpk9uHaNXV
ob+W9gqMu15m1r+Z6BncnBB63yLxducZVV2o+N/1GvtECWBw0fPw3zPEObTX/Otq
J+VxBzYUJLIhuHFyGcPREyjFJ4TXd+D1kVHK7G85geSMe50vS6waoRsXKA/s60J5
nZyQxTKKOOntr03KWQgQN64TakB0tr5/Fz3bsXi8VAfVUE3JOpPATNw6dL1ILuDa
TdJrKWiBg6ZJU4S/EJAqTcctrRl9KFnZtm6HX59amBIb21MJbikMk/+CcsagHcFD
F9NLG6HhIDcjcAy4Xz1NcVmvx2rnFVd2D1wSv0faQw1sIJqyKIQD0NMc4SDQQH7M
BmTFTdngAFC8K2+V7Jba0Iov5xiNpDGEcgVHP7ePvdRGaGhkkO0zF5M+0TkCwxgB
iF88IdbrgdhTDMHBcdkZp8aRvTuC1Tfg8thN5eItYy9LiI73dWkP4ST9dOONZLju
2azivlsj0/G6DYo3GXmrUhxsSm3pi55hsprCXysiBj8GiZfn5qQkqMeoclqfx1lk
t8bdXt31Cv9P4GBSJwp9g3w57sK7E2cnD9FXGM7ZlNk/xzdCUnkHrg/iqjB2EZ3v
N4bZvNYF5nd1CuvJHa2mL/n+NZlMzGa9oSHFJzVEs2n+xqsDtvr3+SGwhOuvjUiT
4128cPB5wbKTsXK5SA8WmO5gFG2fb/Hj6nJzEeZAwk+NCTXIB2tUXy+dTrApW1lr
aCRaW9qaUv+8Mi9lE8hgmcyinDaz13tZ00oVjvloJftswDDWqeLAfobdpZ4TbSvU
PpJWLR1tAy2HGcd3/Mm8xEQoFhQ8os5t9Pu/80aN8Id+JN/0kTq9EQgqFbTZvm0y
3wWKUtv0bqlyL+ls5nPYjC1DrnBr/asVCZkr9z/2KXp8RhJN++9x/Bimxh7cA1tm
+gm4/PYBcpEEFlyEbIk5e0ssq/bq74SEdo+QhiPS4PWIB8zN/7Ugiojb36S8ExVM
vO7NCJP9p0n59uWBQgkrEYtzxK1wJVwfgnM7O4Swh8OktYDUN2u2Y2oSpP+1mlJ8
DZKjtYq74uQxa9Asg5C/z9cCiM9P/kFKO9bRe9LN/d5/VIsMsWyZDmZwTPpr51Rj
VGfaveOyPFcz/ZIKkJ0Tm256S4vEw57bLafrZkRMK80W1O1Vl65Wm7RCTtc+kFm8
7jwtUrguAFFJ7EmB/LTECvYD+m3Up39qzoIaUCKpYmnF0sWOmsgsnbaVQEETcApZ
4N6GZG3Y9Oy8beGUXTWTsIYa3nF118XUs1IFBZG9qTEL3lVdrmNJEjsrRYMhBaO0
Mp35lhAOLH8TVipx7w1uvSaZwGaOd7XM+c0B+gfsjwBNuS5c/6pvg8s/lSPvjLFH
bYdwN0pMcqD79RB199+Tl1ee/LwKw5TYGGntdNl2cAmkaFNpbaKgCmr6glEod8OI
qrsR3edYtTXbhbSBSuo0VB7hqE9MqeeO+fisq9OFsY1+7myxJdvKgXMpiWQUujpQ
XceqlVnS3if0LRARDf2BbG23kWud8yUhj0HZyZCvvj6tMcorpcXFy5FXY4ctn4jn
yOuAOoL5ftG+6eK0dmonW536cVIDMrsfeCja8p+E9R8UGO/eafS6Bzv5cN9EwF11
J3lYsYVGPO2myNFq/nT5DewDAti86TVlhiRsEnCN1ZTXk/cG4jmsljT9yyD6ThCn
6okyX01YkUNHTEXm4lU3LBPMHcWGcliNRaYlMe23RDHo0+EC6dle/hUiP06Golxt
PZLHHuKzcAfUOkkwWhgndwGf4IbECCxVjyqfmCC4ZZZ5NfDMFwJS1IPOm8Oiq+ue
uZ27RuZ/NfB7HCVShWN4xvMtosHrhi3dsprdjJ1iJ6xvwirBzEX3sPdNfix0rTpL
5KvcAcd5cHJl/48Sqr95FPEC1C1Noa+haKE9TNCxVJoJdm28AgQVp/e3jnsVF9Zh
IclAJjZqzJyqqc3EjFT5nJVRklZoLrhpU5+6Z9awsLcW8CP0bRNEytxmaMvAv4tQ
AyugxsKngzo4DYgDgHFZ7I+woWCt/pTLEYLpslOkQWHBfXVpuIY1yPmZW9G1PHLO
fEkZFG4j8HtNpF2p5BlEoh/vgghAKr3GB6SdtnwLvJkRbLGwgHtDMIoKjwE9dars
b6QdydinYqNKwNxrJQ1GzdYEEncUH7BfMr7YfAAeI3S4CVQKbyYrgaHLQUuS7cVu
3bbNop7lNbqNzpSvsRiyk2XjhrPHSulhzde4WvZY1UG5djWCEUR5Rl+NDjkr/WrU
RdCCqGESDjvUI/K3lk8nY/2b3rtKmCcZnVGPxKhbgfqBR28I5diWzhNUtQptg9Ef
XBDphSb2ozxG+k+J195+o9/Dpu+VJ9d6sGZ3ezVrSYPJr1XOiwvHUkzVArbpEiGo
p1NkewG7CjKUuksIyypSxpUhu0gcHZQD5XbXqbalRmP/ElFwh0wqkgn3mydRFROh
sbzDCqBrZM3GncJ1jVhiuzZeIsi1oeN3tFqniWLKmOBgp5J0IvgZjaLMm9wFuYjF
1AXpHswuZg70atZVu91Cx+2pV+FduP/GWiHPOda69EI3F+oL7YggrQuVqt6cT1V6
i9mRENjQMbkNSIK/1bd70q6O5BFh/b1OlpBnNSiKqRqWxC64UETthdcjudeSoj3i
gOUVGpatMKInt+rRMdje61MYgKIotkCWhfXyVDMctBQwhd+RtVDmvo1peZeSKs75
oRUm+dQdlqQM90gRink9WDbD/4ZXMLMR8JTExZEvZp8bcvsIkcHzBUu4LFvm1hTC
s96SGimmPsWw8rO7z3YJxpNzaVwn+j+BeEshfioB6NcyfsqWSaUdSWEevsM5z8HB
yhT9mMK66mYds2+Xj+PAWSoSg7Obi/emu7kdDQBMFo0dMP/s1WB+VUKTgT19puQF
bya1gBReY6JZWFvGxSe+GwmicZqQpk3b/3dviSHvfjHqk9VNT76VP9BsyYPKw00R
ceM0jM26qRbPYttnhg956i+1qzpToHaJp/jXGNaGn0QTE3w/BkljjLVNU7FdB7dE
x0VXL9ah20I23nzspluog1uF4/J6Vpi7s3BFt4jm1pQYcCAt1M6KaooVh7jHWDZ+
+gNIAh9pzCs9xzM4V8R6R9t8kKW0OhtwBQnLEno6Mk3qYXJQDoXpdJ8Xys5SWZiA
m1MQW6SQ2+NEiZNwv3AcUJC+FKezcyYFNKwB2CaN3EGZk6H+yHKwe58+hCqhB8sO
72a5fWlyCNInLG54BNLMrndPKpSPYg+3eZJtcTvsBcrAV34HD4tit7EzhtUbtv+U
i0Hnrf9/sIw0uyfDe6YQO7E+481lRD/1Y1eX7iip3Rq5RHgOZNDa/QvCkGSl/iW1
sIU8vrsyKNK/4lLFdcc5wsONSrMVeqlhuYSZyd0QzwPe5pF9LbXyOxgAPKKJT7JI
wEi90zM78Xk5jOalcmr7Ufpc+sQjztOiEGxs58xEhR3T25b5AVxN/i/UjJa2HwQx
SeJSvqEWCTLNLeTGs53N93alQYmBvYVQ66Cafh8QsMRGHgveAUl9E97UzxhaBUcC
0n17xD4a398jh6wqgDJYSPqylycYYIXbDKJapHewuVMgSX0gxn8/QoIE6WVLY5/Y
j89UGSFI9LDWj7kMCqBA8+qjrzYmKxBOvoc/1v+eFbEqjSVdM2z0Gvm6gxnP6aKo
WAALBEEQtjWxgWQxASXfNri008pzzQtBKUL4K9LJGGTT8CeF6Cv/uZS8LkNUMj3F
Hc6jUTe6QvwMlxUOZgEe2PPFag5vLW+cKbqS0oFx+BY4xI6gQWq2YFR0yFzm2sSD
Meoblu3BMg/xsZK7uRCUf91iOTZ0oq4QrdXxTIhAQameNOiSXVe7GIyjoSGpPdyE
VGiZ/mrYbjSW79mKLkPxyJpW0c1+xT95atpTePHLMS5/7OVwmgdLsD6XD2loA2b+
quUTq24495s3PS7S2EeRAaKx310PHaU1wj4C+xhjVGFVJHnptcEo1h2ZPZogDe/l
iOGbP1n4YmNZeeFcYTibbolvQv5GA0QL0rWCI1su69q20dzaANVabtCFnRD9GyZP
7Agduew72WwxzkMjPUOhEwBmZmjclolqK+Td0bEqt6B08vZnLzJjG/nGeyviXq3V
vwNjsV5mSOHb/ZAYYPipJiUp+MT/VSceNcvK8Tx7x7RhAfFoyCOXpZLpEaLMQRyo
s0loxw0jZq29iNVWcfCeubTNSTIT9znuYnNFGxKTcDHC7zVyrPB7tbDP809Dd0vA
B1dCAY7luUvUK7NT09yUTBPJi6a3dGzeythWjq1savVYbFAW87j2BoduCBYJTKhl
J8OEyGdFEeklQq0aNAOlXVETrbTFbbeXP7tWuqUlLB1DrnoBKpQSSFXjRqbPyVEv
hHY4ps7vj0+jBxkeji3FIodDW51N52czKizBq3XI5Bf4KMgHTEd/blwU+BXSMbYS
qxgw8iinan02XCxwFvllXI8/9xEBV7HhkxG2o0U3mPthNTl0ijfmKlXyNIMfhR+o
6PVcJ9AqTa9vSHW3WYXtCM7dFQTV3nZ3VE1jxSwr/KadEMvblzEYd6G3aL4MYi+S
lyyevnArLlJBIu45s07OjraFgE6J5BMIZ6uBCr7G4KqQ3W4LTfFvVzXSCcrjZLiu
cXv/XJce3o51ylsr3Vt4J4JfkPL33rdc43PE1UV5oRcBxnqKjZ+TiFDngIRnCLMh
JJpeB7JmNiiTu0KpPg3gM7OmXLp1dIOw2Sc3ImC4+06fUO+5wna1LvbmgpsmoxAu
wFAALaXgvvEIP3k6BauK0eet4Gx1OEsaplvzQY9Enfg4gQx7lUWIPglgvdVCqjnY
rD75oT+gDKmt5BCCKJMdhUSfQutn6qnhYazOfY6CmZ/F9b4ouM3IxLljsdnf83Ty
Ug440PZMyAoMxg5THm2xCTa77GMTS2pyZOVU4X+8c+Ah69M3zUfmn/ookk6dFrQ+
gQwILcyKnakLW8pgwn27p0RWafbhg0Z3sMeVePtPpBiOM5X4xUYS6TyJvhLk0+O/
T4G6rUEbiF7CdjPpaxWlSuOd9rkUP1+EuV/8dos4ST3v4MEj6tJjTPmfWGLA6hg9
CQvbMCXnuY3NeqiCGOI9zgJNVCMYsRh5MXc78XvpXb2fGosajRGA6DmsK9Wk33Ke
zF74lMgpVDdcara30jIq8C21kDm99TMMDfiSqEu1xSok12IMjGGcdKwa+W9l+xu5
N2CLidv94Z3GCrXR4wDsmHcu7qSYPGO3HnQaOqkqE+eaDM/EvploU8xmVZo8WMAw
0K14KEpnLAJxxUNhRlu7g8a3EhnLY78X/fvLopoprS0tJB5zLAGElt672HHIJnWU
FLOUFdWST2SuTEZMCKlkOQGt/BSTRxaH1UQYrHEeDdI4eyxF7LS9SZe8P6v0RpgY
hsknvfUfpvvmb0+CFdyXqptNf0XkTeE1u2FOzgQxgKBWlUenVUSq0myL76ct4eER
4WnFuSbaYz9VHPUhbE11iMo3eevCvpneyE+nxpBcxj4+pGA6fHzg5foqG0BTAPtY
BkgZE4x0lG5ofm1Se1IEM2hf5/rT+LsmO0WjMVoApIARx4wxSbbw3W0U8erlq3/w
+Xn+j70dsDndK3GCP9+djnxyXzKoaZe4z/qmJyC4UYNvzJooqEtqcgKFNQGpF60x
Pn8/IGY+aZb09FfDbsfrOJfN7Dvz7dzRFq2sux8wFRHBp2adL4YISL31cuxejiDE
NSCbFDAt0xUrtV6W5cdnBtxR0ll4yZzCB8zZdx5JwWnG4Nyi4XyleI/e9NY3BW05
5XEPrhWJH+1BzceVPd69qhD84zh2Rh7Ni/upnFHkhMobJVd8uevG/o890I3ELuET
yIwSeqF494jBfbHoI7nZ2xz523dXRGWqQBnFUgqxT40iQJbqqsHJ1k1MvRzn4kvU
eCEYPFPG+fSP+MvUqpNLFDc9Bh1VQAbphe9X/UTSdO/X/ZgUETHT/pzd+UhV7tCO
9G0/+DHF9W96tLizTOhFfNxIffWsxGhxidsW6LK7ya8/SATQrWgU++0fb4iOP4+P
uq/G2gNHQ710ri/5oBd2QPJhvt0QLt6yiZFpUmyL+5zbswq41BQ1Ynz/zr+BcCUe
WSJmrgwNTQ1c9o3HgFgLLsjfpzLMj4YqQvWvxzEiZQUeN73t496lZllk8pzk4OQu
i7Ze3RCs2Zfcwu48XhBf/E2dkcWjC9o3B+mWSc16yqHOj80Krp44CQhj46qb8i4b
7LYARDEzkDdRWO6cJt8L6aqo4hGE5heWbWOIE4/eLGJ0b09t3ORgLDAeo7SIDFok
/fJOho2SevlF1V834yYECjauxqyRdLl9ErGFUuxLIIPn+Y9RpsRY8QMKj7ibw4Vt
2Zh/JSlJ9VTu4ml9zKdYAce6PA2LSUL5UdiZL7P4E/LgN6j+TXpyVy4RZDKhn0Qp
zlwK4RKsCYCHT+uuLA13Mq7WeUN/sI5SzOeRNFUnE06zzplyHI7lHOrvw9kNTKSY
nIG9qMdnyWeYNqX2l3POKBB9y6xKJhtV0a/3WmpZLKg+tGcvTIoSQ+u9hClyooWS
8EVlgQ4LTrhU4IcwMFjkkdjfA4XVUwlSYW6rRlaqdyg6AK7XB5sxj/2/UJDFCcWJ
PpaTu8TPvzXcS8guoSSPQ3Ci2TdvUUvo4LcUCllGa24vgy1EH9Y3mToD36p/rvTO
oOfSlLLVcFGR1Gi+m9hhLp9ND3MPTSM5IbnsFRYEvodMgD10V1ZDt7Y9oi0IEvX+
/puAt9618ubXfzp6vJ3jcQDxf9+4NvE6P2fOItKCvS8aqxg4dykuhq2riztLzsWu
st5aaQHBlXmuJYqzGtMBblss1ZTPxWdgEsXnqDiWtny+gdx0+AKw8S6zu8kogk5y
LeBNzq9/1SX36aJiWTpKXy3Guv1R6o4sAZ8+cWc/3GnC01uaS3wc1gGIHFFLasih
IcKYHk5l32LmVi1/IRtCF0DbZK277NWIcjxzCxGpewDwpzDhgnZom8Am+hBA9+Lp
UpxIVmu4QsIdumiz1ezIhniIWS1TJpRxA7CtHiXq861habGPPlbDyj+fbaLTlf8C
7ktukSC9kyxi3cGE+I99w6Ml5oKYpNVQqULYJwd3AMQq4BFl4iGNFf1RhanSlFEQ
ZxqYGO4tcGQhI2WMufbxvT5XztbhDo+YLEgHaaO574IO/pDriCDPYn6XF5/Cn67E
xYRiIZ7IrF+y/DmSwu/2OimPLZQGGTHDtZaco8t+oc27GDQGhrfMpM842QVbQ7wZ
9CkN4HndvrBo7KS6kpYthkGMXCr6TrNNjBldSjXqqCWrm12/JyX8wP4j8YmxrzUV
tcLAemu/XFM9GFdPHjgKcEVqhJrcMz4skKi3CTgqHdGIaJ8WwUsEWw1jbrHKg5Cy
7vUzwEHoLAw/z8CADqLZkGVDbqerme/eXx1Iou3vCCvDPqpQZiTwwysA3IwBk267
mCgOUZsErdg6/her6aEOJZMYE57RL1EoD+wp9rL3nX1t9h3Ydq2A2uvGdRAz+W14
u5xjyD8Vv4d1ekFOFsJewu+u845ojpAQ6Nj3oE9C3ZkxAcHSXlKBlc7fW7twwicR
joqEavdWa9VeOLLT88WWYB8RjJAA7k2Ubm81KlmbvNqRqTC1pqdFmy11G+F5xMYF
G7xbFRIwWR3m49unzC6eo0fCTeM6XPg8UpFVs2C4P0tEO402uriyd1KKMXqPje2X
Z8KlKYeqik0OL+dfLAjLjoqWW4OUlt4gO8dzBhCAV/xkho/lNgVOXINbtsMjb/0m
oszIRaxb8dRG905NKTya/47BPZOI/46QqZwRwM9pfo6t8QGJQuZ/JpQNuO6pC5yI
T+agvV8JjI6kQ7OaLLtmZan+iLgOqULiO9sg3xqXlERcxsh7aUFEb3Ei7OW1nJyF
bqXPWaqluo/WCHcN2fEHA5+4aAXbvn5Tir6scI5jmJ453SnNOpU8Q0oAR2Gbgdn5
z0HwJk/BmYgOddvjkL6NxuZ1hrMBvuPs7wGWFekjsyNuxn/gDlXAnBq0PFnvFqkY
nwhWHl7t/LRSQX/ydtFpjIhzlfa9IklOChfbY8KLRGconXFNXFtqEEmzjiak7rAt
ENMHpMFEjyOD+fJq3qlO+YMFogdc1PR69tFfG9TbJQBqwPSAvtMu/HP2Y/jI0phx
vGqM4Ga4iHSWzTN+EA+wn3QEsfIOWwjQeiYR1uJMICmuVVkkekK8FbKD3pnJg4ZT
aXc4WmpS6YziMEDa+4XYEFo9AacoUft/TAemz5cLHs2mQXjMkD8J5Cpl1FN9bgHe
VvoWHt++SXsAT0+x4mpfzMjXtrQmNgFWgBP4r3HA3NETblOOnvbaKj4amVl7Kavd
55hG2WbaPcyARg1NpD7Bj7OGXn1vWIWzs9MHBMIe2FTg9y8didmOfX2uTl9aqj2X
zL3wdw8XaraQvagfilL5qs1BQeTT5n7048Balj3zQD/hzXwAIbAvyEdfjKED2CO2
qpw4mn8wfFM/7gdWl/sHhAsfhxLIRG3CBm3b6QhREnA6uFrD2Q8bkLGFY6q0fk86
e9f81CHduJ7rsNylnXUeTdrqEetCJaIrJ5VV0vY3RgEORxg3OnTRIC/EJ7q+WBN3
2FN4JBLQJEpOSpzuDm9vLK6qggsMaP/w5eZZm0l6NS+JGGLN1ztIeWwuk8ki5jkK
WP1/9mAeqBmmwPoGurWRviJYlq/vhFk1X7SLxC+tKK5T+TwOa6+meaaO/4cok6nA
6FCeUQjGPXTPyisIO6xfg2BA2B1nrc/kOmL8LAlAY1V7x2do1ykJW8moWkbrA/Yg
QvT8sTfE5LB6bKGmx23tlMa0ipIKTjRNZobrYUEi52HIVqtihmGtkQDpnMHgl2T3
YmxT2ZQ/3Gda/HRRdavUo8QUzl+T0E1ShwNNrcdxSM/Txq9o+eZxjFChgC51BZwT
HpL937JuAog6C4fQPR7jxbSgsrl0slr/KnRJqN/3zxHGWLId0x9lnxoVIYI+SmHJ
QgQCRXY+cervxQNEfe+AmuB32ccyyMjzbfFZJcxOE8gXTic6QEn+Fu3CavFziWfR
DXwTuTfthqfvK9pCKfFF34p2tCxtzQWllW4mbXbFTTHXsTdi0omLpkm524LmsAFn
nUjCbQ24iFfdKHo/s4JAJm2i393u/L00mSM8SoGri2uzVXs+eTIem9S/BNRtNsY4
0s2mfwCW9HYZCMwivCI2H/BWvUI0PgGuiPvQ0b36FzOeqXrB1PC6V2f6VO+Q1fqX
qnwzX2i+Jq/Vj2kTzt0BN0MW+c/Zbq44EfK8fy7cnW8Bp5FMknJF1t7p89iNt4EG
Bz6De1uR6a6iXSBwP2P5yPkN2BgbHO6sdRpLBJW4XXRWJZmaQKQ5lYIoarwT6X+U
cXeKvpNRSB9XeXqfuekVPlD9t/Ii8Miw8ZgSRl+RZnk7YC0P7ks0gpbQquj+Yxqz
zhpHLKwB1WwPgY3earLAZuDaboQRChtJfaAQHEs6/gAfawYAsMJy0UCWrg6B2DnM
SJmTeLz5J6Cgv3eK1XOpNK2RV1+SZAszlFc8z98QKKV81KTs3fYGYxBiY1M0z1sE
DlAkoRf7MHsroBldSYR0N/eNRWOEcKGBY17jMzqNwTRr3hWaEyxNG+v5hWYzkH9q
mtigyr3Y+IfAvte3/OOoLbro7+5Njk2HYynu+rTQusvxePzFnWFrn+UZHR0C114D
RCabbN5ivYb28LMP0pmjYncTMiTVTr+KzxKXD0+Bd1mBZonXHT8p3uBYoU8jeLNP
n5M6OyYlxKnKJK2/h1gW92KBrwPl9KVwOqBDfuoByYZjXRDoESK865z5TOilj5T7
kwTBX0CRiZxBNZZZW1dOBSvLDeRmXP8tzP7FSjLbTdCEMrq7Q3+qDvoncSLks8M0
GcyxVautOtbbKI6pY26RnGCv5MdFcqMwIQpfeymyWOTl64+7l4PJBxy4mGVY+4ne
uUq0d0tn/TaeTQ3vs1m/BsnM/NxsJ5/podd4IDmuBTSpcC3saHhLAz3Bhmxme48v
8+im1hNraOnHCp62CYToxuxqwGfJlUjPS6VK+maZFTFgyrvXPYWkCLtTF1q0pAFV
a0TIv8A6p7wRzfK+YbKxohIYu+2O3B2p4d9lL0s5/D+vhxkRIdcdqHRVgX9/ioFL
HftjEsRjGqwEFtsuCkwzY5gKCZCE0nBUHOQ09Xi4yixo1b0uWWhe9aUmDDJLHzHT
QbNNVH7uzYLkp4ebdKSvBxGrf6Nf6L5mBXPI6WFmuQKWHC5SnX9g7wAt/PRNrc22
yCIW0bawHXh4eFNymerlBkcCV5O0ZRwXkYQFihhYZMcx8jkQw/Yv8XgcnW52FzL+
4/oW0HiMA3GLwgWRxK1UOC2xoscF01Oj1HGjS0YIbFKvotmk+bI8fzfIDYsv0J/u
DvU5Fr/wX0A43nca1/5IXTHIqT5S2ZAarkvPMOIE4jMWUpe/xHgjmMgKVCA+PpV3
eWAb+Bazcpnq8q8RFEVNj3fa15YcYgMFohLGGn1RPa2LNDw1KRyOWGVApbqC1HDO
oxOHTan/cG0xZ2GPYUdwgO8W+f9ctQ0RpLjsnIJMo1eqSfvVxFk6uc/7q8UAlEou
9iMXAQq7OuqPRTy0LA2CZ9cNrkJWmt0E6MKKPRVqCFwZ2k1X6vc7c+60veMa6taM
rlXJqWLYYqMiJfgEzb+NAB0LGOxoLJ/U4RUp9FLkJ1Ro3j2AAieZGx8expE1vV+t
TKU/Q0ddeQ/6Yxwns1bx1S7Eojqw3wqk8hHPey/jy7kYUYKpNRfjaCeb85yn6yK8
N6PBED1vPVIQQZrNVJVC8BsurO2RiTIsRfzPOZlASxfJB7kzK8UvTCuNf9JBt+Qv
XBH7wMgt2/n4GKYGAl3w8NuroZbTwe7se/w4Z83igGGhYTCbzrIE0M+B/RsqiK84
IfMCJb266uhgfJnZMs7XoZLD6vJPzUsWVybA6dapayZ/e/BcjPiSOYTGkRYOJ+F9
0Jhoqsg78sJWImaNfImAQGnflr0yhJTTuTJTre+4EnslkUXYLIqoCnM5JCmkNBJj
7xlK4imeOL9kdGXTfD2l48gELI9p3Y74G7718QkYk/9tzcM6J9GOH+olzgq7Hw9r
yfOV5m0KQsQY0t8l3cU/xYuPlySrgbBhF1BnJJZyXw2pQ7JMWhw6KjTRR5/vTRyO
nTBq4O24l4oy4x+3kIgUdbWklmefd4Fcn6x6NfHDCaIrmX8/4ZnU8CMGyBhdqxUr
jqLV5q69BjdLEH5HKvi88eeMyO5v9fgXrLE7fXTT3GkMI1OK1vKzz3n4u6Cm1TIR
8HupnPxDBZvJSzRKvxirEnpk63PP2R2HuwqrR+b5VkFfYkbZJeh0Nhk85S6MFSS4
wMcBLA77yXszeMJpz1qC24q2yQqXUcHOjPRScSrInCGYhut2XD2rq01tMogdQFX0
/CidC/OVTkBCUdzFMCHzZ4Qcq/VCZm1k/7kYjtpvFdA3tsIzOWXZgx4cJap5V3kZ
tNV6biRyfh6zbwGyZi+A//xNNql5PQamK5t3KX0rTxfyB8OcKjAbrpQtgIHSKjUU
kLcZ2GKjmvE23SlraqhuVoKPfidaNBS0i8ccx+XhokpT8gksEYMeHAC5PYQowEg2
j7a8lDRm67DrnqiuY9PtOM1rC0Ow7jpg/FQvGixUJNHOdO8DgAsFRBdt0beYNIX7
VbKbr180/fIDLy+LL8eP9FfFTxsRp2wxroDiOPScTdAjdlX5pAFfH+csl4WRLnqw
K4NarX/070PD6nScqeWrTeVriX8oOMc8x/n9m2Vp6cmV22jbqfCC97M+CxaceUCy
EgHlz0yeQBBmLxTuIfRs+hOZHpqmA50ZPbvpwcy0duvv1UpXlHrIQhpIDL337GXe
+Wmgb4Jh0zfzXxF0WSrgFJJLGKKQu5HPf5bt0+ckiIV7UqIL04HwXAeBLL6EvD2r
BQUEItcTOd9auxp66sw3J1t7PXUFOwq2NJpdxYNY5vSOGFWieICvjc1poq+NB3Sg
x5yABMpLiFsd+BKdwBLmkNGvecdcnuyPES3bfhsWcOTAm9dbyNjXjEin+0h2GPb/
Kzyr4foReUFs67PCgGhkPxBbTnhr4W0Hbbc86125si5LPaLK2jK7wuFCuIO1Oue8
1modqxsIKeHZTV62jmKQap90TOko2VL5DxIyOAv+0YKoRE9nO0W0SGhBNUMkWcYb
F2hbuGxqud1veFjyir7X3TEkFvxaZN4+wHTPuQuclHXOmGdN9B1cJtW/rwO493SL
+RQyoa5JzWSNHoJq+ckjkoOYf2I1SruTeLVehuA08xECVIUWhRA5sknQ7tmvyH3E
8QKUJ7VtlsnFcxbauvL8k9LC9Um14MWlkMDGBYi1HMTgYOek71OPhvA7fzj63hdJ
NdehYc2TX8mnOxyxRfHtCJEOTuGroi47aik0TmFdBFTTuyx9UeAgXnlyG2V0eWku
guXOGPbIRWSu8vQJ1GydUINDE6ths8CB7zmsz86Ej0Boqu4x0OiO2483p97rrqN4
XlxC8p9CY2N1Sp37ifLMFacCuMB56MYmVPiiLRBN/FFKzGv4FGBGNgECAW1mu0sw
iC5eoWSxMm03aerFD7ZuQ16PiYnoFy0TDzh0M7KK945WUCIhHJK6KT6uORwXKUkP
uOol/8Md12fyEQchM12hPmBPNBInBtPdkub9JUDrn4wu8lb63geUoZM0yGYz7PwW
lTkCZq0K1Ml1Gwe6DhKQjzl8Kk3YvKux2LikF2ribHlFxa3huD5A49PMsqagmo0b
NFxgBLBTUKE8QHLfC6MsFcU51Jgk+hLdg4Me77UngGJ1ulvHtunYKXgrs31XGIOC
qwb56f7F7WcDBjtAPaQ5cPWv2D9JYhB5b4UyaBnsGMWvgKzZUAi53xUFfA22AFbQ
R1l6+kB6HD+xZkkcZtcaFRfVuhVAqJIYLYaxzsSIS/VLcUgBgVpocvcf6HQQRzdU
wSyeh+HOIhg0+7ijw+TsPgHyXfUJ99J8/6UIuB2hIl0WUO7QDP5iEtb9QQbCaPkB
xf+CZBagkKy/6VtL7fKkn9aVkltJxIa9coDP+mDjVyGwzCbKVRa07NDyjdNWyfu9
D5QLZiaqJiKp2VQ5ci/h6DkXioRkQUEIxoUyqoU7kIxa9eIH2FXfvWbZCEeoqOZy
JHCoDomHcLx/vw5Xn3i5ya/uapSKhR0RKnnTwjRWQFVp6Wdlg2ZEZiX1zwND5k96
MOIye647WAtKevmkqrNPEqB81uwyMCxQhwkP6MIq+IC4SQyiJKAIQRFqvOu7C3Hu
gNH78flo7ErpevXpkCJpEn/9kH37g6+i7qh6HEzHCl9ABuOyuvenQgEeJuZgQtO+
SsTwh6zuzBXct9gdahEQnqOefm9U+dBCNgzwn1HAIaR9tfZuA1ANnm7LVQLHViiM
tDG3fpxXGLS1AfvC6NJX1j0PRPLZeIrItwnUKpp0LLY4U82Coll4th3b6vrWemlz
OzLxuj08OW7AGzrnAfVpOJahksoH05iF1xCWkmhoqvRlQkoW/XrrTLQyPersnJ5i
w4cunRg9juxVFQuOPXk67AvMaOtfO+y5sAcNCAvK95jmpMwaVsY1HH0Ync+6frKT
NzbeUzgyTLIdGWE+6udWt2poZYMTE+6utTXRGg4DvYcE1wdZ4mDtOOedmXDJ99Mz
cRpPp0506tOiN/CVGlVhW656ZfxNJmdl6DWQDtHSHI4K3DoBxowBcCtfs0GG71jm
IrbN4Z2NJWsfHxp/Go/ykXTf8DNbRJXTgSImbPz0bc0QtByZ1go+bX4AoPQHR2XT
vM29PyVa85AAMZI9i6vSGhoQfMfuToMtr9Z4CUKJaEwobmtjnNzNnkZ6E0Ltq3hk
wvZ55zRlvS/3QxEkkhz8qzIRrIvzWwqtWPZQyA15XO10tIhjSaY9nn3eJCF/qRSD
SR0iaLBBCLrO4vAajB6LZwGd9Rgc5BHvFlPJGYzirc3cSzLlkFK8s2sVEvu77i/g
lKgE4G2QsKIeRAJpesrPYvI4456rYyfrSTqJS6gmTnQjcN0yC1bUwZ30aUOz2YBv
azC4G8WNEhBYyOg435nwl+X68Qhf2jHORrVeq2I55sJeMhJBDy78s35cldDiAgqJ
ucBLvy9Y8jJx+suS8IrYVs092dnJNHhKEFSTH5Ay5Mg1gVzCBcCwO4p1xdaLDuiu
42J3QR2e+yQXDZIH/0ZW+3ZXqn0Pt8++mlpTtuQlnI6jXxap9xlegU7HgFYCBH34
glieHqb92+8QNa1/DqCZnkIHDLvlr6kTr4sl35nszGYyPURD5DvCOxGzJ5I+/NYs
x1DpJvDjnfJkqi/v0et/OX3qls6Z9R3VE5mIqRRxzhGQi+TPm9inDf9z+09mpvHj
oJbtGXsGuO/CgAsX3zhU3aEo6EmATT3/aVb42/uXyO7KZgb8rUi+CTcfPxq3wloS
MC0ifG2eW2rTAyI58vmci3bE72aK1DhADyKHNT2yeJ/54x7Gg/cL25T67Nwuu1jo
mfbb496t3A2X3Vnp/cobTrwT2dzTkC0YZ7HGi0P19eCo1+fIxoFWLyjwNaMx3tGu
izoBcePhT/zd7BFFJmE5kOCe/08MUtQonjtHt+cT2cYMPewxQhGKMwBS+Rk+5DtY
Iq/xD+HttvzcL6JRQp61M35UtjxpbIJupcula6zFExRk/x42x3g2m3EOFL/wJDUe
6t4TtLeQWHqOa/NGsIqYzAuvHRj6OC4YHJBFngXmYQ4iZkDBrWN2hBVN3hEVN84U
vvj6HyrYDf+Ju4+qYdpVNLSYfmo0/aqTOk0zbDxvZqaYl7/zCrPUXYXRPR9ocjhY
42PPZ+iTp2S5VXFGwG6hImS4si9S9ADgBqdkbaYUlqU319/u+1EvadVovtMKTgJx
hUITz2b6TC/w67HWzgH+EMWZwnIXiZD39e6xfxNqIbiOwgLHACB+WQ5dkwkrIdHo
kkIIz2bSSPz/0uaZDNKJFaiH8G6D1CoLyVTsP86f4I0N+h4jhvPL1EWYPT4gpV+1
w1i9cpwtr/1wO0FU+lRgewGeY+ql/KJZ0WJCVcDGEHyiM4+ogYRJ1tGqiLcdUxqR
q8HAS8rzzt0UOq4X5+e2dyklRDeDGUwYR9Q/LP/CtBqNIEpryw6qNRbz7sI+38/U
I5PcblNzfgLXXNfqncM4BMSlfaKm+32Iz1KNTzyqRUxX32Rwqb953jsHiudkOUkX
iPCSE0qoXTMpTFFkGNdn4V0r5i2xRpnPMEZtAXAG7vHeFKFk4NWjl/LvUnpyM/Tq
aZlC8rX1NsDoa/WGd6BoIm/f5EtOwyJhlKaMDoRGNmPfBS1cSsEv0NFVFbx4beEz
dD/5gJmG98NMHFMs95PIOzVNv71uOi7zTTbWTT/ytBR+4GfaQGmyg5fODCQ9TrBk
FXwGoMXkw8NGiiGj8A7W1TZ8xXYR1+HOHnv4pQw/yGbVIrpuw1gHNcGWd6xxDhSY
S4SO42+aH6QtoD5WOUkFS2hQ8bkVNPqj9o0XCtd8y1QokIN+onRSgP9I0MYxzSgk
WD0ev4qPCgyxCaDFpdigyOkYAq7dIzB0n7nMIMGiIiDqHGFLrtDQegru3aH9RE6V
ow2kgm+taeIH5QDZ8j+gwzIV8LexQ1c+0syU2wVkMV3m0ZMPAK8vkuiAoH1OZMWp
iKSx2GcjqMcTRu2mylH2V6eE7flD7Ld4bVS/ipNZccMnN3EzJGCIhbdHw1TvPnGi
7Gt+JAWSvXtopw5h8eAqG9r43+Lo9AhEESJ5oPn+ZPu6HJLOLrOx/jTL27q4hWFm
yXcFp9RKCeH7qmCwtzn7a0TxyCbTkFls8q2rcjP8dIxqGqJYPHaKe+VP7kRIAK1q
4u1QTvsAgyXI0Hw2vWqYJG0lsJrQQbb0IX/f6DujRAsmEF/9qvHLGqCcAF7Whdc5
1e99ie1dacK50oV0RL0bHWhAsRIGKlsSvgYcX2sUwIoD/YK/t10lIVspvZW96you
wg5irnPuBxnBPZ23us2qsiEMBFw4lkh2GwTAoRpRbsLHKswDBq/l78NOcaJxFeww
nD7h32gG0nXw+6sRIPqh8V8SZqbiRtxd2KMImuabLSDHzI11Z2XJEwag0RxxXJ6j
sWmaHheNHo8kisvzo5oL7f8Qzt7+j+n1mZg3w6ZAkFLjCcDcXMciEQjxWSr7viMY
6C414oAK7i4LQs1VVn2IvYbzGMr9Jd5u6rTcPoAM1qvGtBkxoJjMr3Em7n/PikLU
rTbB1ZybBUT85oaatg0+3pq4+hOH2/c9rVqdMwG+XWcgN+00wMBZyBiBtamFJK0h
pGKwCcNkmqD1Ln8/JjVixsaxvX6HdR4k5yOg/B/Pgwbqv992DGESQC4T0ZEgvObQ
Q8TOeVkhjBYT9GBvEBx4/FejHkuC601VTPKPCCVR6wqDFyUTbrHYNGJ/uAx+pHE6
xo/iOCijGUmFmAwEyNMwaJnCsaGTz5VPVwkBZfVvJr7bm3Sb5jHyytng86OKUcet
g6Js0ONXFE8n7UbvlkWBCZlLkmgB1MU8tQMEuhI4ev7/aLysSAPHWq9LR8pYsQ2s
YxQEmLgG2b2Bd8JPFjBN838w+Ho1vIA4HxiX6uHauYWEVgXi+qVT0+7d2t/pD4vv
S/Y0jUh/SUkxy9UXn967dyJzlNnqEko86F6rKje8VcObL+6vy/R6yu+Ru5HVFhdp
lnLN0eo77G0xhDwgwtwaxdEb/RwyHndfqcKlEHTIDvgGzF51ea0C63jQ0i3sqpwy
eL07jNdf1W2a8XouiDHVZRQpVw8GS6ioJNtQ9yT2DZTdPBaaW4RxHSgmH82zbRYg
JRY1UgoLWjJvJ1ztrDYY1IIYRYIOryjtlf+IP9HOnDJh0nsKqU9L0WPZpk22MLss
nNLGrjloq2n6MdPFUx7lVAIzg+/2Bnpq931/ex423FkZCuQryrqSUmZQ91XfTJMR
+fyCq0a/yoOZWru1y7daMehRfZcE9NfzFeQ3bf1+FcDhvwsl5cjRHoL+wwPPwTaX
pf3tMWMirHumbr1T2FGY/mFRSeB5QhrRwKWLlkWJmEv8/GNQOxeF/0tMQ8RB+xoU
fU6YFgg76abU9NioapGaHO6Oh7FjD86X7HwIM9sT4sC+YbG0uGPXv/JccMqRuf08
EWSFwJ+/bEOIfgKRtF1gXZTqrD/mI+CA9/sTICN4/7uDR/P6p6SxCaXxRDy+tvt8
izg6zywpKoLRpEcbX09yxTe0Q0JT7J4+zNzc7bMpuVn3uOPNs/4mOpLXW/gG8YuT
/vuGREUFI7XymI0rh6HgMSDfoewKp2hcxTYPHPKav/t8fyAki5mLAyeGoJpw1KMP
tXNd2MmK2HiYdXDFAIgdp4M/IPz6C15SJOiZQovSPSf6yaFB8J8PMLIhHzroPqma
MC1s+f5rtP43U3pmrbd/kde5KF5zWIYcPLLLgyBSaqdmjOW4SUOnw4DkOQy599fX
9DJtWEPvpyCMsYPttSBrIV/AFt0XWW45nsHc5OFAMEYhlj4TfUCKfZq6ZdGQFq3/
w4hA9cXAFCs+xPNefdk2doFuQLdWLqc1Fl8ILduUbrCBJ2C5AwAqFo+8FV8wdr9v
FzNbp29dUIak/pqCKMK0lPnzQqeqWy+lXOVlNHfi+vE3ttAsiQvvrYMlW4pXXRxB
Nzbg43ggKWCd/3PdZq1fpPg6sTwVSgPRHAW4ohc5dJ6j21v/IwpEI0C6t+CRN26/
7aXyWGcOxMb/Ezs/P4y3Q/RoTjX0500VQ/RTJGqtx15A4SakLECCK4HXQxpTlrXn
wgqJsfq41Yg8U+WddBwtYhF65bnsdq8kU1ws78wtmABGGbnShwcZFLHrF7KuWG3K
EYRh+rizKnfV0Q6/hgfDzUgzaBauXm3CRYSHik82QdMuxBcewGtPoIXEZzg0C5s5
Uqqe/EaO9UGuBEi0E4OVNtllzz2PB7BM2YNKqi1zAQkW5y8237neQOhsa01Xk2a9
znuUcKcSuHDwV2iVjHyg/2KqfdVJcW/rFvJY1M1CIzgKIPfzZJSO8SQQI5HoizTz
MEETKXAQw32shdrAqpXabeeMZaezSkiY5dFIhz3DxS3x6z34yGDShIMdrtj2+Z8H
Bh90Pbcd2xCZbUjnZrp4afZcvbdNtqVO6SqwBlytbKlt4UnqR0hrL7scmufURx7x
jhpF/GLl+QDhvFmQUqSym8P8Z0ZpjZUieOttMx0G8QErodnxA9lkSbAo+9PBmTKH
QEPCyUKUPt4wRAUuEbCTSDh7ocYLGrTkMZFsN0PrqTji5qAw0hlCWbdLw19nSvPs
FO6flwbqrQ+J6G9d5wPIu9sF415+Cyqna/k+kjizpQQ0e/Oe9U8l/KKzzxyT0JlU
qvUw3OGSwNu1Fp69aR+rKMbz8h/2GuYy5YhBVRliSB9kWTvNgNpqEGAyzxGDru2S
2xkNBKZd9bv/8052MJO+bHAR4RtEcM3VEwol7CCGRcXc+uiQAWfKlSPX5lmAwjmT
IbHmLhyo7GRwYwyVSA3Q2KkezJ20TyfbQ+iko+5euUay7yB50IwyV2/OagqVMye/
m2+VjdsnweHS8m9lBXw6/3mAnddsq5YaRIWpocRikJIHTSTcLACZ8/hfPtgtSk49
Gwe2S65iNvLhecyopNFi+5PSsEWZjOSLWLy/Sa4irqpncZFGLG70gRq3DQ2ag6Uf
IfFfC7AU8qANEUMgw6oF3Fm1dV6eVzTIUBINhlisRc30etyI3sDzCGo7H6lQbtAv
fuJ+WkblbCbdc8kjZDEkHXXucd2SvORBrLCWHZLmh3UGgySTVLIoqD9/Bm4Vbn/H
V+GLozfbKV2Nuo/w23az2BOEvpxTCQIz1i6W+ofd3MMVSD4vhEOHegjSvxwuTBA3
/KtpPnCUaLMwdocrLpvcmurLX0eHRjVhjExSDZOkx9ytLmXHXYNoNyEhwVNUKxzn
8bwRevhLXSSB6r7MMvja+SR+jUPHvEY5sF/0PFfwVYLLvOlgDl0V6+OLS0ziWp5z
TgWBlZgwkbGDR96jvEFNtSJ+xqmP1sm/aZg0rcX3HiDGMheNcpTKZxg99UamS/vp
AiqnCS4Ir9uHe6qqzVmL00/d3G5gSesUVkmxVBFbz4PtzPsUvPmqKC2/Tb7yX133
4O/r7D8V1V653HRRE4t8nJFXuzWo/XfO8jCd7HgolNMwqG+S0MWxte1clt1oCpdW
YT0ImAkxfpwG36vcUPL7Za6LWapzR//Nn+qNhhJFEFAnjei+VA5jy6Jw6QOCxcVe
rJOiuevunYOeADzA9Pi8tjIztbJpoA12KDhu7lW8exGxOsgT11ytDAWsYgVoYZzP
Xcn+LsZUlGrjHc2sntBxYYjBJ0waB23fuyF4Ret8yFGtk5zwAR6GDT9vUa3u3Wg/
atqCNmu7uxt8FE+kosJfAP/ci2MiYYCfbCgCJcC42o+8alljT8W/LTmkrDTJZfq1
LUEh/lp41Y5C4rw6MbEhTuGj7zuZg2jJsIYsDlvA1SspVQNCq3E7W6UI1NJS1z4F
ajOQdhLoHYP2KiniDcJ1OEVDeyRDEwraTdQN/fk7OrYs8rspRUCCCBfMHs2ITiQl
cHOysAyjp1vSqLumlggypZQCEP1ptkN1r9q5W1uOdIJPoLuadVT6UQCzHHPa3mFK
mCzNsNkWrvmgwQyRx+YCQFFIYlDb681IPxukws0h+nq6aWxQAN9Nkb6HyXUpcXxX
VL40v8FZ8mDURFyZXZcxR+PnBab2U6FG3hswy6dTnV83hQv3vzC+eVfCSiAi4Tn+
KbfbWICV2+JoFX1nzUIhlVbvR9ea2ALdkpxoKi9w9lu/PlsEsOeDYoC8xDytIaIU
0PvfjA2K1XQtVRG6ovL3RMknFjZaU57th7ErwQ+khaFHbCkcqVHTtGvGyR34JWdc
BhxVvQwq/AWUjZyYUN2gvhbDmEmzt6ZmQvKaVDz5Uid0AmLnKWK711cG4w8t7OtF
276Vw9t8zp1TId/zZB8pa4H0S4bO7b+w4dnaPDVoqNv3ATEYXS2MzvO8Us+0+bDK
RFYq2RlIuIwh1zhCvVZWh0N6HmHy5bKS0u+jDtPpz2AncV2zfsXJ4YoMxtWShT/c
+1q8q7prZeSiTENpAWOBIGoysXNBmn8ErmXU8f8n7WCUm6qTv4+h44HLxTJtPSjJ
r+9FBGczPfXyAf8ceA1/cZ/kbgnJhJqnm1BLHYfe5V4ZKm8wH0uJnvK4M6cQm56p
vlv/UoO6733LqI30IdRDy1u7h4vik6RhYrf5tdXlshOqqEXKLnivq47Y68APFKQA
UgOlKEaLHWaDC954FzX1/yCgs7h03BDi6mdd5yRbjoapWskAtFCLnuxL+LGvAl1p
L1eSsvo3hIM1B/SVQUr4nIQxodSkaneOciC0LX1n1HI4BIGWBXMM9nVHfTbbL7iz
SutoNNFv6rU4BA/oV8UNGninNpYbm8nALKzerxyblSTDMzkyg/NVpaOcFx7yvSp2
KDuABD82A1UdA/AnsOrVfvXVhCoWkiwhFBdc/ZebxQa24y5ouRY4D3BnoCYaA9cb
m+MFa29zBKrSGcy4DT08zuGi5o7oHCImVrOMU6dtNqU1Ql+2Se7BXf9ZxTLBgcjn
OXJi/zqMi2VFTPfIWnAhdLExQfu7PutBlPsdTYfqPUMxZGKUH3isB46qKqCL5iJR
cCK2EIaI5mf33ijgbj8JH1NUBsU87StBoP1BJFkY7HtKeIG7ta3vCKaKRXCZL2od
vkFS0smV9tonjkHsrb5HAGtSwURREzDX8a2uhmubprfto//hroyc29Q+lFk3RP3f
Amm1eroRxa+6yrm9vb6bPBsFyh/C/RWpbsNpQgJ47Nn9kpkbK8VFu+6cgV6XpBoM
P61nVnF/c8Ut/ECn5+xiu1jKlzmGYqoxKW8IElyCHMi8nzRyZsAV60v0vgpyEAYk
eaox1Qfbkgnc4IT9ZguCYUYVl8/9Hl3/GcXQIk2Eni5lxlqq7GUHv9rgPxZvecko
XhrgGs3Blix22+UTwAx/qPrKjDnJ3fFBP1r+I3W9p+m+YweGkIpoJvdnETD6Bovr
c1E1Vk+uE6J4Q6Fp/o3sQ70J8YK+S93m6hgW/XGeWYrXvnO/4DfXpJQuJrbjpzcF
NMinZtvq3Ct0hdYi8jBcUTwpcrgfVg5lOAvYQZaJZBpObqnWlxHTwrTchzAYtW6N
AZmyXHP07XX2MWCAULHTd4OEb8YN9aGIPYFK4z+hz+fXwjx8rgM9VsfPlinhPUvn
72YjqsY6su+lzZmrLcHqa7IXA9cuY0da6BGAa+4zwwoa9ILo9n1GNBk55yGc73L6
4oB5ylEguFvFG9msQtj0BReyv4qbMZUJaSRuXk6Gf52dOLXW5HjapYqQ9iqdpIHT
WXuHzc8ZWaZLSYXmknwEzH7NMEtflQqkeCoAQMSuqYT5LfDgCUhBjfmsZXJHRglD
n8WbRohZTRH60BVBSuSNF+PDAEFsWGsoNBCTlvfSXHmE8KvWTFmD9i7BBJJwlcJf
mpggPAAjp629gAcp1l1uL+uysQ1qlOMMHrapPTrMbNRNVfQ89bg0+nwaJ+LrEVj9
+ojNIPY8Isr+EPV9npl73AnScFu3QZYwq6TWYQLkz4cLZk+QGPrv/IdfFHAngdHh
yRZI/ne9Ywvb6qHg7GTDjVz0X6zpawL8vdnUyIvsqiXPz0k8LC5Dc0en2TM5Nqsp
jqySPdP8TZAnoFtRc3gWiKl1eoH0SeuFkCPebRtXGCg7mDvQ6j/G427IZ6SR+yNC
9BOWNE+oGyEGXB2heETOAaeoxv6fXCabeoik5jguBpPD3CktibdW7EI4Xj/qsFLX
/hteG8A3h7KQD+vpKxFDTdOT7n8HOy1J1stExPzAqpw8a1lXr0Sh3aLD8l/f8xNL
T9B4i3LotBvzq7ZmU2/IjCtT84RPaedQ/0KuMUuCpdvgQgzlvWh/LTEhb74P/jPh
1eqJ89XH1GN6ZUedHl/cpSxIQ6Uil42Bt27Y96594Ahp6l0E1gU7AnpPTbg0gpXp
rIZiydQ0aeYtl7ZJANeo/a7Lxmmkw6JZE+bEc+kYTL2NaiuHw6C8ncn+k9dAXuaM
3ccUCn1AtbNsFrb/SaDRWCaUoNZLpFS/Ke12nnT0P8eJNsrVoor/L/8t3GxOQkYp
uDiPpA84Uv2WtA49i/dDmx5VqSRxvoC0PQPtpvYrHWQ5u+OD3ph+hehKR1k+E2aN
u8hl7MzCeZNTHTk+TPlcLvd8DLKKrtbcIOyBuLdBktrUAHiqfIcNl2RJHvfTMGZx
8pg4BseZ0SBMMDxCDvOT3S3L6BE1uoxQb3jhr7uRMC5rcvik5E2gqKyR9E3FFGoi
Hfqkj72nP+/CKiiSoKR/pe2QukIO2RN/1LOXAIJPVmXFyNr3QHQ9yjayUDp2Iswy
87+SuMvTn97xtAvhEByV7JAygf9mHqCnxrNbIJ9b9z1tOrJY8rrSVmq4ONFX+ZeW
GQjKwzWduB7TvhXako/B7tIutbLAI4A1VAfiJfdcxSOtcjmn6dPNVx9CGGsBh2ES
a0WbEOaeNxuYu8ioJeeal5uKY4SDDa8Z/XSTqLsKlWFrl+8d724qNkV1l0d85E05
piGnxNg+cIy+6fKXI1emwiUdZwic0WmfUVTB1/z8W9xtRlHUNUdGLqzgV1ZS8Sk2
n4zbrOHDEDTCY3ergBhWyuQzy7eiwGLzPKBY8h+/WIhpYR9khUtxq9KtIOZ9KHtC
UkyUQMDMghBWTOX2gqjYoXJ6+UuK1TZV4LKwQLQnVFJWV4MKVl4M1M6LsD9NL/mP
Jc9YR1FsqNvTyHGBq/7hYy09oyAgzapkadcAcvYqBVZlOwrZ7xiVY/w3CbceHz9f
z8XF+H7RWDTv2cz3PH6Tr3xrlBqsoqcV89NOkJh/vt4baTO6evXIlAbCBYBltbM0
pX0YZP6zG1Ej9YfVTKSj2FSrUq88Y246Wx4+GKZ1ZASrDjr/cp287lvQsRevGTWW
KTuiraEJNUXUrLP7Vihfy3wNGtESF8DtAI39n/7GfweIGyyRUr39AxQfGwHjxJb5
HqFT1G0a2gzPpmWexVytPccAZgowEXQIVUuTPBgzzbJ4VftKW0Rq2SCb2Tf1iR8h
o1HqcnT0dO1j9Tr/N+n2vsNep24gChCltitIWqJuG9g5c6ZbymwYjoy67VmH6ouH
v3S4fmq3YcZDcQ2mihI2apa9OJnujajAl1qK+eLHzvsPsiWx9dTVfDkzngzILyrC
UNUnNY6M1FIaY3cWBNzZxKUdIBtuDSM4rQH3yuCU9dxEJQRqOovwg35eobZXeRim
J/JWHqwDzvXhc9baMh43VHei1A3BQDlJG92KymoE9NXp7Cs3A9KEoIjuXfuSMJ+Z
FefDhxAnd9/zTIYIpwS5ow7DgvmxyTNru3oKw2dDIkY8AuLS1q3It7Ke0ow2QrOR
A31uGTwlLwLZ1lyijDGdJMPuMBVu6tjJONWLDBiszb1tdNQvk2qF7DwMarBFCv9e
mfyu1N9r1sTdPCO8ytQjhl/PrkoEHdVzDKzDN7KjKfc+n5TYq2GWAJediZF7LJIV
hC8WpQgtG8kMxF1Ov1Eys6jGOcksgXBnsYaBK8h7dr8ACoxkX1UIlDdsQN9JmD4y
gWYHiE8V8kke5vbSOr6WR4FD7yqsw63g2r72rImozPcfyMwOfpYnz/v3XONW/0eM
E+11iiB5LyEKPGkLGanVWHLoiZx+NPuxKl1OFIxb7z+kh7M/nmAa4+70v806JRsv
y2YDkrqfY7qaBr6bl0Qod8cFoaJiNAI+ryzS/jCESn7JXdUewZg1XQJOtC1UfjZm
Mx/027IDHsHUxm0ca1fj2ogXJ0vz0Zcu5xvRDfM27yR9Xv0K+XISc0cdasgYfIGz
j0KAUnA9w2TnjZG5Yo7Gp72IEoho7yE6DF0UoFhNSGJrDo6q83Ti6hB4cYqWVbMB
HhjV0kCSJ3UuG+nW1X23g3ZGvXMGtwIZnIYr8lEZLxbN5oyw3AnyLrwY3WrqF5QI
K52TXppqwDIKFJCZ0/FmHRoiD01HlUL1GNs9mrWtYTJcNJweJPuCw7az9jLvgYDi
pnCNLLcQ90zKoOtXI0y5AT14R2IcnQILQDhE+ppmtgn8QGiMGr0+sHXmc/3Sfmrn
vOziKTgEvfp5wlb42p9+SJyoYvoXCFw/HLay4G/0lClFz0qF4wy+k0aWW7tw+kJP
I6ThHO7/PjOfApheR1hMYUsKi/Nn4U2QN0YLYDmGbPCCRy8mxjcyoQIiF+PrLkpc
Xq6OEVDWd1HHZZbqo0123KtGcJnSM0LOeDTHPKEv6cjq91R/vvwzw6Iftos+X4fl
4KRRScnM8PoRWjoccot+FdusFcBNPnT7p9sw5P31FKIOoB8N+Rpq8pmeYBIwwHoI
HfW6ZrfRtaV45gk8iLMju+PHeLJ+oPiUKp67AlR+0AFXaGohwPnUC+zU1bJV8/5G
Zfk1ukLGN4F1CMkIzYYYNJSwIr52AVgF0mmfTrwf76CkdRmQzb4wOjgKa8rAgGOI
ExeFELA289LkBdE2oFcogjIfzltwXIoVhE+nWoSktpVKM8O5rvhwCNupQxwcpzQm
Jd26YYz0nnyuovsHRdcMxqrfu4rqdajajfHxJzOkvjQn7mI3oJun+fmsC8jQ4Uca
ENTK7uRK+Q6ALvOnfeQmtQ3pzln4CHNYtejOLJby+tFGZZo5bcKY5LMqhbBk0bmb
xZmZj3KSbjiqq7dSM6dW40nBlFydm09tx91qC9tpsxveWHT4UTyNY+Kn2DjO7ZgQ
FzjlAc4FVNyEsDLXvJ8HtBTJ8b3fmwp7ZLcc9ZmX7/awKy2ewazOOFbRpGZDKxq9
D5Y7KEut0dY8BhA1VmX5OxW4tMUqhdUF7pilHBZdZjnG2CX950lUi77UIgULrCPU
AKbYQyNGny5vP7lSYZHTifILCvzv1E8eGPyMIXZ6X+WJpClbUqssiFGElsM6MWxF
CbyxZBMX6SQEov7togXsxDvReV0JY1SN4vuwtTc1K1xS0GQ4YGHl6S53TD7AUohr
zczWjHo/Bxwy2jDOJV8jxcab43uE1D1EeM5asHz9geqnfXglEazy1xAMSep3QaML
8N2CxMhMzSL9E0TnEPsyZF6Ak/YOy5v5AV1Fl0KatXaqhr2soAGJ27KLkvD4e+MO
r7J35H+TnjOa+cG0+3f/JQXZq1mm5G8XAu6haj/mjETrUPhhfkcrFuLx1ddNwQcO
qtC5oo3FALsEeeGjc7BaIQrlyrJ0+cBRA5MJ0TP7tCqS4X9+PzTLtkxMO55+OHV7
vtEaOEtyahS8ktUpEG6KYPm8J3O3Gd75dCznxprgX0mCF4PusE1a3Ic/gPHtOjHq
L+xGHUoGsgUfY87j8RjD6YD3wwgDnak1gLlxUZnxRhBLGiXCPrurDAhSxGZD39cj
3JxHE3P/RipbaZjgs2gr+H0Bc0sKHEg8k2qlTrnWvRVk/3zHgOzBRb7hiiK/aTGu
x+AL4PmKYwtqUtQwJeJGcWcVVrz3OtGQrrDY1LXx4k74V8gOaKRgd5yCsazeGDmG
dupCCm2psipPxszb1zLs8/c2hSBpZb71VI9o1VDmIdnMxpR1cmGpIljx0iiOj3Ys
lxQ3Crpsz3MkwFTTPn3/NzEOodVMvO2cElhUSdfkUBaghQgSDyNZFznOwKL0c6KI
8po6uh6L4Zm8yzqhTovUbRgEaVDnmi54k3tuZ1wRRJOcOnaav4vopGpokpKF/tX7
hsVLnOvUBi4sVDel7ZHzwy4d625tneGaD2C6FVVuHNs2QTH/R5BfdNINtFDImJFH
burPVBCcLRitWYkQB38zf8eWe1lRCHFPvw0UMHXUmY34BaswbG0gn62qTNR15l/o
juGjpwbk8H/Gh2B0IhpN+OucSxbybiYdnE5hJXeMROZZXxzcn0gnztfeSytW6ZGq
KAR4rDI/5vBICxD78onLMYX7ZUSe7W0zQ3+twg/3cKiEQOiQQfItoh8hl6bWFa4r
IHN/NuEJs7ax8/gKbXA59Yf3DuDZLs435nNykdEHhi4WSFOvIYVIfas1rLDfvfP2
Rd1Th9Cwx2PFYG2CFzwEAxL8ngg31zgyO1p/7sdSJ71c23GJC4fEsTZ2xTbiRI0D
lTM9Bfrw+pzTweVZ5gzlnNEgICWboqu8TgfTXwgYjq/nIdPDYV3N5ugtxT//bF9t
XoF7VpGwazT/3RPcDNYKwA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
F1fGZmTlfSAPxO8tY/XQNXLzgg40H/RR7qL0HyYBUa+BoppT9Uc9B8aPIf+wqlaV
ic7PxuYIgXMJmewZW6qv3vigxLG/L/TI3JtxltYxsURDh7CP8MN1/Qeu2M/8gn/3
nLXIpydKwe3mgbrpbqshckHTl8NJ5v2pxPWJxWUn9JwufWaImWeEKOdIJZ6P67p2
wCiEZ9MTmUZec0rrgqarEC4RjmWa83Kg21vPai8wzlKvd9lqusnaIC1SNZEwSnUA
B5rl1WssKJ95QwZGPr0wkMpeGamR1r78MvIA63b5jGvOlPh50sjXOTgLB3loujap
v2qTHXgtTd22Tj+eS5OKtg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 24720 )
`pragma protect data_block
brVGN4WbUtyiP8as2hlKpdIKlPF+9m0xtpbvszQqjTmo3TcZfL4ohuhffjUm4Gr6
qUYJFZxQEo3Htc7Xp79UhN2eSF+VI76+qqX/oNdLQ7n13o5L/9SoRvHm5bEZQx04
9n5vTkAA+RPWMePau+X0bxeQH0RCXdOjZcfOQTRIVVXQ+zQUWYHo4GRF/qIZUqCp
YJi9ZZIrAs9+jteodyg0OOG0ywFeW6Fm7hZiT+a+yLfTcamnqrbHz6oSijwM+jAt
ur+uS3iBlp4dBaM3rTs0GKT9a84mf2PxbKRZXYVQQ+WjQhfqckHrnz1CZl8v9J7o
JAk5UbWu5oZZaUM1zldJEn8x4cwmx/uO08UH78NUJx9GUa9rdsTvSe5AHNce4fSE
v36IQ1ryYs9gzKkvg8kR/F542shYJppLK/9V3quFJwHCnVgrpGHfcerpsMIrNTyc
s3zo2raX0Wjvr6H82Fgrw/FyHG8aAOfq3omdFp+6QqyGkToLtPLJinOOXKmhuzcL
58rbojTd1fqGHYWyZbCrMjMvMBzRNNLnpI+s4XZZbc1+9Zmh529sdD59pLNMfmH+
UYNBi/dLOq1y+GuwUJKI6yNXISq66tTuFbc4KWLub0QXrwXX6RznHHdsyAn5PX+k
/GfwLHQvSeliqYExbF4zetTqPdG9xl8PdssRGA9ApzEcEwC1UOCr+/zZAlrZCE6Y
F5UFEJfgdm44Wxr+huMg/mvRu3Yt5hUcYvFO5XR0SF1XR06+wXg7Z+mexGgsBpA/
xXsQsYrA2ElKwLBYcvVEy0uajPfkhyN0Cy0ZBHxqWU1YxUzzF9AJbzhu/zRWHWJr
g3gT9SDtT5HZRmFqsSZ8V/v5z8nOIX5FLYPVtV3VMfZvzA+PNn7bWeNIfTy33wo5
FkZN5Mjcq+KAt3jW6WRFIJ1zMqjkJtnPxbFENaR2mxk2FheYVfvFCf7BcQ7YqUdF
YaMjCG8x0Q5ruXGzpP9l4kwUzGiG20ISXzXuzBVw9zyMyQ1v0zCbeM8qNGbZTv9e
tGZcm+qLBPfU5B7d7zovHBGgosAv4MFQf3QeVfOfE9QmGqnj53LFy7ngWzrTHc1p
Ja6KtbS1qU1EwooeZ56N9fvXeakc+GU4+O9EPlSSQP4Vx7HMjKaskrkyjhlkIuNA
Dd5vWaKzTgYHn9BOVyiN6+9HadCOdTws0sMkgSFPzjGXf1cviYUva7B++XCDcAph
hcXaVid7enECBnuBF0gaXNwqpOnpm1+gvok5II8Yk71LC2vDzV4v9IUBwFQdTpN4
/NHOwcbzRNeEgQdqpJyx6m6vMhI6OL4xT30OnpbGb4KJH9+xM+8CenrVrQc5CNxp
Lm2xFs7ZuKmJFPpChk0SEqRFW/ml0dMvH9vZhlrPHYqqzgwqZ7DaLODGMQXOk7xd
nmN7e7MacNK6KdJBilNpUMFgL4qQ8YvYfhn0KVnpu3PQEdRX222HCLqIx1fUmbV4
YYOP6HGoA8vPAApYIgi9JLYQeeam+srru7O/Gj0pDbgq1rckcn5lWF19B5G+cGOI
+LVJPMxIPjSkBfthqApLR4q8scy25AqcoQUqExgFvPSzFD8+CcCbl8A+xa0QLsmf
1sZ7rEslRDRuJ1j3qNA+gfad0gKQoWEmuJcpDHaQcySdcZmbhQZAn3CX0MpIZu4y
L6NSfNC6HMBr8K0w01mUzAxjUOY/9DIW4qtVPQ8QnI5lxJlhOEu24MK2TzqpAGWm
JmR1xYiGqg5cqS4Z8bc7qZX1qu060S1DdPnb3TZdxyuykQHDfjzwakL00Jjig+vN
Ud9FJa9Fms5mPkZvKQl9lfRyS3JT0/IBpzj74Ss8JRE5Vzfx/A6g3Vits1hkUljG
QMTojfpT7GLmVrLcWuMKhWjQ+2ekpBJbEbMn49FguNn79xQTRjLlth3EHYHhh5nL
EtBBOYJo4JgN8YArjVEamDGDBE70zgY7CZjacuKwWMt9ewCh7ibP2JWOMzpBryf2
X4Zu8/Td/YHd7QWr8z2RmDpUJpmErT46GJ0O6NtkgeSwCTkLZEmULWYQ1KSuQlvK
m+EA0z7pMnXyEt5/0Anr4AW2JKuFIJr1I50yvvNOICFhuMACjqmqYa073QZHn0So
qNKB+esjpg5jE2tZ6GT9fTUh2G89oDFb3ZtOlReKOVvZBuWZBhiRlg+Z2xPP848g
Q1f9CcV0XqBZU19bizgQvRrRqSrJ/EfT6JhSzOhXtSG9wO28mRrYeYWbONsmoeGa
d/KJ5ddpHdFDIRTfOUmPE2DJdKzwwp6SRN8rVOCnFfh8wqjLq06SxyRLDJJWWOct
dR1SNHy1cO98iFXI7LN6s7FHsGYjQGSRCpXWSj76B9wmQcuAEF+vCEdTQlLQEqO1
T5A2SNE1MqqEVcbvLpjCqFS5VAPHLTZkSc1k7g2U0yC543TyF5DkuDlO9xZlZNUC
jrqKXC0KO68Rx2grvEDrPtRvDfG5YuEZGMH6P0h4wHA7iWkW4iJa1zqqqvo2M0uR
rhoSNfZGRvSSMu6T39hkzH/65FKlbOWMe9gLIUEM5bo/qiVGboXLaHPDrzIook/1
os37X44ZnQ9TxPDFkKpifC9ONYrnnSBoNlThS0B2Mb5EOMo2BwpKKzJNXXpIq1Ed
IB391u9RlYU5Ee494g2B/Z6rlMrBOPFxegVIu47tIc63kHFQ9DUzK+/Ee8jQuV5J
lNfRPjBOZ9MBm3Pdkjb1R0oXernI+e1D5rEFvZ1R+ogjugViSYjAQuYqV6BdpzSO
3ysTeoU8mS8fADHl4A7jdLXsvGH6UrpYYiXbfXpCsj+/7CTbh8tpUrMWUrkLenbR
jkNfOzimU3hFJycmxY+zaGNF8lyHJqgWUjqIengAIqq4ai2jB2KjdWstuLJNmULq
BrVXIFrj48IhwHAoTuQA/YYbcsRrNdM/gofA99lQOSL0r6CvgT396UDNWDnKD7Kn
PLuxOqU9UJFo4qHcK8VtXbDibT6SFz7Y+SvVUj4xXgEKyhn7Hx8KVfL5tEuynIp5
MkspAu6CL7uWpHMvXkbHd/pyejcUUbxoN6zBk0LU8dLK/L4sDqoqzGj25onmYZVb
AnCvK0gG8lkTTeAJQJ/sSiU6ksGvp4eZmx9HG8UkwZuIwnbbpZoUTkAciIT90RoF
81XySS3RKwYBZoECyAje+HNI80deUUpuNsg0hfWcI4Eryk5gnK5RRINDX7Gb9sCv
djVc3gHDTw/L6rXzeQpxgJa+Bra2Ahm2WSKJaoxJ5T7910MFBpvmCLFB3I41en1k
QxoWXDXTVpJlyvpdd6Te+WyU3xMIlk2hkXsGI96R0rl0/UWracADtNTGiME6jpww
T3bgHTTc+lDGUt43bIh/JbIUcMw3Z6oa1iIwLD2iDrGHLlcdSAw1lm3biQOufMSi
OM5SlDuGGF3d7xz1ihd8i5Ffk6sEx70hU70c/t7LHRRw5CnlO5XajNGeTjAJV7rK
sJpRp9iYS3NSpKNlW6lo0EDOYAaNZO4RaPQIk1y3iEBXbVIPMiIwvFEJOX7lN58J
UABPF3/c1M6yPxUrNXtttC+l3Ws+aAY9X13MSeLgWfd+0Tjj+YFn9GGZwoQkoWWC
TM0TTtyQkGwPVeyjqFdxX15H4Ut35jt3hwWfJFelzw3ujuJ1WoARr0w8p/SL9t1L
ya9vxFd26zbQpu4dhiJRbh6ut2lNpeWfuvtt1WfZBlr694NiPoYqwuMCnr2peKaP
SAME026kL2vKl5OonvZALUWNxpbPRf5HbgRtJxdz7Vf1ltCtVqm7czFkBUcvsEKX
/cUXq2QKQnuwtZizGMPPlj9jEGcOItUiyFWD/MtKGNOi/yltofgqrtbnd8CZ3jPs
AcbeqLlzPtfHiDRSe2qu5HsbEHKrJBvaKtoZK9EHZkQGRQbNMHfWfMRwdtTUP357
PNR2283sszt+Lyx6y4J1WlQCABmY5C09qgFq3+aAz6NJMjytxaG2EYKS/vFSXJc9
xzOY2EIQvKWE1hq4GO/h8Wf5ZLuu1LZmjDqVP+1KHXtcXdhfjPvmYC5ku6gZ7+K5
JPmOVb/p53Qctm9Q8+x6a7N7tn6JY/M6orektxk4W8GkQVrIqjfV4Kkllqj84v1b
nsWigGcQYz21ReQQqUKo68xm7DGy0ngcRzKlLfFaIKK77cmNS8GQ0fEpFbkl12zS
xaHXdt24BqX3XxxvM5BwH9EzNBU3X57vyZxQxNl/JE15bZJuLgsWyx4Vo4u4GHSx
PX3OVh5S4kXNE7MMZEQZAo/9Blhc1S/HjZDF+BizWnLBs2oeDp9EpJkHzzgpXVX7
/8LZXS4DAJGMd6J3hUy8mkJVmPr3Trp0UmJzg1N5SvSUe+32gCr4h7Ac4fYdlKIF
4h0hGwOWoJnTXsvJWqY95JOugd7YRbly9BnvS7NmtrhDQ4A4Zdh4fbE4jeQ4OhNr
he72L5ITWn2XXQAdriyiE5IO96rHrZJ1n+HQAgmV6V8SS9jc1Z1ojnxxh25Fs81l
4HoJ2W6OWZFVnFMpGfz0ChAsp8BnXZgpG76tgoyxvxyZMrRfs1ym+YvHG4r1KAtf
rVm2kC3DqLoZPg88GBU0WSqXvvMH1UGSQ/OHMBTF6pLEj+B9OmBFx/8tNOOxJezG
/LkmV5gxqnOhxa7kbghK22dPR8ocSzoJ3R9UudvyxOK1Ao0+wSHfC4RA3BoknOPP
cz+3diqhK25UlxgpoWh0lHw77yUzO4t5O70/K50XOaOdFCGm39vBovDAONP+dVGf
oWKBuZwP4Z9lq/sD/If0sdW7n/BV286vhGaPfEcTbcS3KVVzgDqTePovZUccCSsd
NlxZVVTz2EL0yJy0oChKHsbDX8Tru2TfJLRU0wJhMaeBNU7HzEYtSyYqVAuWIdQ2
pLDHMWzjr4zZVh6dLy5kng4EoB/WnGruRV1jauaxBKJ51Hut4Ut547a6QdHYad4l
s07HaMg2wmwejABo/zNEZk7yA2pGl/axrcB7rUSzqQdTbh5nMIDH42kruCcHquo/
pagaf2LFEBdSrWgXxZhMk9ZlIDQAO8uMOY5b5VechWptznF7r/S9gbcI+5v56AkO
SigiTPu6rTfshcFmntaD3d0dB0Ir6znGb4vai/KCdlzAkak8OtRJm8ZUVjTUYvKe
7xFinrOnZrk5FtwhebWyDYwlYZ34Uhs3I7PMF54yVP+dJk/pvQZQBVlKkgtmK/gA
sBBrlyFQH0FiWYw/nuSXB2o++VUcr0KXxGYmv7+UnUBdI7rz9Qd46yLzSbCUfNpH
7F0O+mOMsm15uaQXwawTlt7lHs7T1IjBa3UMyA+NAoSZuk3I0bU4QRhAlFVkjyX1
k1gGLWp/iLDkX+CDUZMGMh74KyA5m4uFHSi0WX46bHtiJutlkmLXf6THMkrbb/RD
Qx5SvbpsSMSA9MwqUH6l1cqstIlgaaW8XxBgdEHhiFwEtA4GE/Oe81rQ2jCeAGae
WkzhU5qRRjY7/nQ6vRpEEutM99m/c1ROqLu6nQ/lb51lPFAX/Gusb7hZpBa5gtau
izkL5A8fR/+5ExAuL0zQY3Eaxaw1IiFyLEOr39CTT/Ckp3S+gZ6dYzV9GelNTp5k
zmZXXPSqOyxB3nWaP5hBIAEJBRKc4J/dO8kscj6OLdhlqxlCbZG8tygDgvwz7Wr5
X/e0cC7XbAGy+rzfiwp7T2ii7NPQGBuXDon9K67odqWjqtQJrxwGL7SrZVBCCjoc
KIN8tRFXOCmSrF2Wc2Iz+eW6Zx4kz+oQVPMWAATo/NX1YMjbXk8kMGWsiXewKAC8
+q3OgQvJTLgAF9BbF2Nngf5ZbivMMc5A1Ce9Tz+qmDXqxiMKGR78Dp0nGhXV2Q70
bRRP72aFTE5yi94OXNyuxiyWEZEHwPbQt8X5RsX7qAYdutA/fAvXE7qvfJ4NtwWy
NMQySlPiKXeteYVxNDGuKw42xF87l9Q1uikkHW1XYzWFvLKVXME92MwaTLnHdBpa
xioKEeJAeZQu3vJr0CaDLxZaYBTXl907jXFI6e+GDN2inCpV3ASJle/4xDD9i/mP
jqEQ0LA/+19qjUzNjEA3kL7Tdkw+B9vflTklmVuXv1C3EBGzS7D+O0ATkT7RU+qb
6yo6UfnGNvWffLUBdSMECaWojFaefeWVd75bGNHsvfQyEXHP168Cmi6dvdIWWkbr
C0FtOulz/ix7a57ljg6BgJPIu+e9IpCs10LnjDjSipMQAkGYroqF0BowWa7H7box
51cxtPqpBg4LMashv9jz1YJF6wt1V2UoDisSqftAttToPE4k7y7kXyIbEeGec7x1
4kQR31OHsousrBlbq02dvETTEh8rK4ofDONg+6uJnGI5BHVR8ZpygH0YOKYGOcIg
QLKWgupevzZ2JJKKShivz0+IALrN/iD29iD6sUHkC/uAY3ZhYi5ujxp7yU2g/DIg
ekCjBL3NtrceTMbQEZXV5bns96Bqg8PW1h0b1jl9fSm+L1NWZ14rfJQPTLD/hubI
puZsHWa3MMkNnKAOg3Cmks5i2YI4zTmyze1Wx+DxVVxAxNbEc/wpUibMVzTaVC5c
PMiLws5l7TsfYQ4ZOALkMrS5ZGQVygMhqxBFHIrR6iEcrKZJXdJqvQ+GVxluIF2A
KpAdNqVrsoT5K4RhhxKQ/ve9CxA4ALkBBqumgXjMtxNQ6m1rDqwb3vv3aZcsXc4/
+UYaAdVlrXzGAbHQk3eD+ECI3cfn2waYKg2ENoJvv+YL7i3nTkzvnjtnLGxmFlcC
+Ng3BTOoSsgHHse79Mk65M+jy9c6AhAnaLBGtQDQq2bzaBVbU52USubAjAPvPd/S
e6NX+h2rvTgjg8aGPGZxRq+cvPLJNAcExfgjczzjzh0iAkhdSAD+jmLZ6k/eLioi
7HFtjyzQrUN4aSpxfiq/GLkrOSCQit/VwULrYJ6TvEGGWCafQSRoq88+WIqI7zGK
bdysLCY0o37biJfrdMOUgC+NPe7yCsZ9VpLtO2ad+wkAHTGSFAxTAB6qx98tNf3s
lSI6Y/MtnHG+wOeCW6ayp9NrhYvWwwdVpWdX3RQw1R/TepQWju++Yp2oQ5LmbIMX
fWDbp2EcW6/XgZ/FOmw/2mouzEcWiWYR/dmViI2nNPER8UeuV2XSf+WVDrrK3dzz
/kQS022sEGLLc9dV8bHdNdJSJAwXP0/YX7CyTVuLOfl+Ll6Ry3oKf8LXMKS5KlxU
y9IAg1dn/kAAEbgm+oSw7ZIDW/SZykJxpIO13XNxEgEKLP0oZVsDaHlDAu8o3yvr
L7ggtPBfipKv1ZPXT8sJ5LlSWAVckrJ5P0UecW7iNLzYQEU9mzxXV7eVVBjPjUvy
TVdGZOt9Xch1oondqyPAHRswxNvJYsn6yDyvPgyLwPlXSRaIvGTcbDa/eys1W8co
AbyvUmjfR0TjYijq6kwslzDGJlYbyx7VrTaKi2mHteMsY3teUrc2FdGX/7AW3tdk
y87M0wWfOBlmStWLGxTVHAqWzQNRHF5Dll3n+6yGaZHMtNKCY5M0daCrS6KaYmVL
zWpkyHyUAeOzyIYWaFDTARuU7IiyhawUxLnK2geLhcKo4uqBeafMqm+yG63pE0fq
a4i4ZomavaPRkDATvB2g5CZiRdA3PK1LG7DZPaN36BJM6RZa6QxhsY4bKDJuI0Ac
Q8ViITytoqTgTAHRh3Oo34NivkhObeWEkQ6ZG17lGPlB13w165CkyPv8IhFK+c//
Ma0XR5P1sXuPi09i9+z8aQeIDk4hLnpK2OVlR9f2CtseIBUOGUq/KF4A18v7mgbb
yHVhfQ46gTX1+m1fZph5cL83dpADySnDLJHnmjOQkG1CT+s7zv6du65VA/nWfL6I
XkWqGMALcowj24DD18SDdm9/SWCwfBYzARpvtDD6it4SsPl/FdkQMtSOpP2Bn2m3
b/m+wEVCjVZ/3WV6K4Gc8ZP9rOlkMtvT0v39gMpu1IU35BNQihkpQydUm6xtBQ0v
IN2svnjAXX0QUhtEG5O7Lw92j14LwOBtWMIY7RwB9c17JdzQyYx8ye7RxBziVOtP
aeyJ9XIVfwVws9J5ZK+hMLvt0Jk8fhvUB25M7Ss+APY/TBakB+B4O6m9j2BBT/tg
+T9Qe27P1HDdZN5hivwFVgAUrlpgMAExcch5Qsq3dE/Wt/J6SeV7r8IIm44OaQEL
NdIUfd6UN9s0h+oQtkg0Wc0ZvmtWfLxfbASBQ3aoDreFTAUADM1bz1k5aSEGXxVp
ofdx0M/lkda4OWVw7TwEFHwXQ+P+IcRharo0nHv04tvO5auNTcPLz6nJDnfBt6hZ
ReaXCsn38xXyomYoRr+J6YC9bMMJNgT7hEnnA/O7aak69dIpwjw3rC3L7UH11etl
DXPw61+9klPBZUYy8JHuxqdIJ1rEoo4F2rkLnwiedGqXtZtJv/MtUnATQohyrfPi
z+1nALANeTwIMgc3DLCstyXxL2b6XJUhZ/ZjU7IIpZopbt35Y8mcdWyBLFGuEtbW
uhZ7rg6uJ/9wCHkgbfZcbhyebxM+KzhG6apx0OLjjgw/ZVfkAGwTg1iYE7hY9a0X
vqbqf0noj0ifNNJ9rjxxsDrCbsqjndp+RUAQTathCFbT72Lkyl2uhzPMKB9WVCHM
0IjaMqtnJwvU2qavjYb4zIboW9VpI4ZZbjHpA91toLK07X64VncFaHP3a5pNGVOB
VLlaNCNaFeuWc/Z7dTueTq14aboZg4gnBrFJJNdeXOTJlvpy5otsZNlvTUGIaEHF
na29SaGWnuCPptb96uawGSk1XAnZPVUR4L8ltc62TCYYe7BxJtDPXQtHaPJmJ0nF
shyaKlmvF3ygKGFRnxaWpICWnKb6hUgE61uuZj8y81tYhIgqwLQMrFVztQjDVzDa
asw3al3R+UYAP/n8027oKSDoydyk0vPUN7be4Y47QXzNtrErI9gwWSGt6Fpnhvjm
0BMjQoJ2yBWlopUXk1T197tT1z7OgeKYT11svj0WeIkFE/2EHI9e6QkW0FHXHJDp
mJnhvBCDG7Ti8E1q74dnTyd4P52bi8N91vz5jkEQ0izh4MR597kVAUfS4eGqJZVK
i3Hg8dSyJuzvj/L1Dl+eXhrrxej9rv5dtFRAxZufrg7WXF9Wfuz7x4LKlf0+S0X3
KKX+Spfuxe/iiAkUUfCD+aFHAlkyOH/XiVPVr3dWNHwT3R9Q6WVIfQMOX0O9J9W8
Tmu+Vh7RVYpDWu2p2qNimYUxcavQvDiJoq9enSM4gIkh8xhosFxGFUss9dn2K8cV
hNK2ncN4fLf/sHhzIE8U/sDXo0mb1Y+2QcUQliATqKZpGJO7GWaTCdU1gWjPviHE
QYjaXy/j8UXE+Ag6Y9akrvixq3z5wl2Ntu0JEekLXHTFXDr2R1ONH/G2ftF9U8oB
VhsDQyS8x0BS4QRiJxOgc8Cpsy7maRI5INrhQV6+MlAZM5T/Ypffsd8hejT7dYC1
PTf9S5mJTTCXE4oGkmLw8Y17mlMkUk7T2EDtJA1C9K1H40mBYY2vcMxI7aezeaQK
504nZJjE0Fui2IcFOdp2iS4qJW5XTsdcMEY90jjy7RS/FsspwJLXWobNEioWz2Pc
ksEFyCqMpGKFlldlSI+D6B0BOMYWZcq0vTwslHYSdq/MVSN/vs1Y0SLebSIHZNpk
YrpBntTGDdQIcOosD045quu8pSyUGaE/gKKmRXNYrjUXJUSSHg0b+xrvXgEQPG1n
nSX83lL5ARVge3Gf3XJh0ThdrQrPDrmQnmZZkKQmjgyaJddigcMycJtm/xuUBRrl
XgDdOHKmth7OfCH/4o1gEnCSa8CPOy1tHOySornR2kv81NhrM1KvInFkx1YUSl6G
r9FtMUMbIO0mR46jkjoNcL/2tXFnWJKQrZT4EEUU0bzxPpxUUXi1a3h8fLU0MQ67
NZVHX8+00oTx5ZEgHJYcHSHIqAH1XuJTBec3g0+ICLcoSLsAUqNjShM8Cjwq3qgD
nXXzIPnlJERNDPxHxwcPgafF7MS4Ju8NmBhhZWHLOn7nzwW8OXtSRqWnFdgRnli5
glnGb/LGZXL6tbr6Cwk5lfGb3bwoebXYuY9UMfZIkTu/UspOBsjQ+BhoOsLdU9Tq
4gDebtkOzttgisNmg4GVH9nfITaMnTeCyGfvYDVjQ0lJWDln6I6r24he0Zmxt2PI
UwQkks9wG5joSURcocMl/lcDUyobG87wxya9Ct9YNJnoL0d/lUp4iwfxivyoNiZ3
4xXfAzpxpxIY/WlGKvsFoj60xcdxxRFCT49197+DhgAn+jvmKyuWrdYnzCuDJWCC
Au4d+f7bBXoar7QgUW/j7CEoIvqPefZdK1i04nr+UL1M+EVnttD6nNfNbyzahLqY
EzmHr+345HBndOP4YqP+xhZ5z3u0tdBePBlxFcmoJS+cdtDg2Gn9Bd91j6Wv3gwr
ojQVxc9JAYTqWbfU9XrcPRCOA/uzzJISA8LXoQoqzeVUecZfefG0flcZazwYYWjz
y1K7pFSLpke3jwN5cgMzRA9pz/5STdSfJIgnBcYjbBRutD2e9z5oCdPmYNhMKSvJ
P18Vl22ugN0639LzHk44o8usCZNO/Y2jOzDT2auYxMjPKIGe5xjGzJxOk7gJa/+b
ckPDvkpoz68dJzgPV72FrAuF59MkFxPruUt3FWGjgtYTqZw62X5gtpHYvda7eurR
BEBT/arNbERUt1E5N8ZzOh0CyXLmLhzP1GjmdN0DJ82/4bHHtre0uwpns26m8BwR
Khs1Kpp1RcRWUKaO937vO+d4mwSKAfCjpPT3zhCxAhUiFlIKU24Ax/uZfwsC+qhE
IoGFsMFeqw8pSfs67nZZNB63B4/sDRjbgc9nbOFEvOtuaMyF1FRHuuNRptL67kZO
918Yy8fBfcUiXVS13b8+2w3NRBVVprXsmBKs9yhJd8UK0fk0n2oQwfOAlG3E6JEM
YUgv9dfl168HtgCIrWPCOUE6avlr4iaQe8J68AfvqyNJr/76criZl9lrWlA4UQpi
GwJmCjNnN/uQKCCqYs6+FgupnARu4jUTgXP14ES5w0V1+5LnTzFcEmDguef4+7wE
lltxbsKJTBqIp0u2SNZadUdBMN3vDmf4O00BbPeUPC/X4j0FmSmnk1O4moCTXWnb
3v6a/iNxumLHjzFQ9ek9GFJW7n0BuWZGImJazEjl4NJ5+2lcGpt24ZKpVVC48f1H
O9Z2pHUnjnLkZtC9RsZnAxgdjQSYOboGwpF1WmzwSgVhoIQZaS6RQbf42enMTLff
ZHpmM5Bt+WWfj0DPbahdAfTxjMPvKZghubZwmjTyMwsPHwhXLTtXpgXUIC0CM+Ss
h5pQktEAZnR7lj2TpoN2Dww3sGLCKONYMK7+5KtkVDbiSfBC8pQMdLXJbZBZfxJQ
J0f4r9NUTdP6TuG6i/YrPyqZiofwVOwX0iNW9lAUSHYbvKM9IoFbFwnSzCX25D0r
X/Y8PYYzxnRBePcnqZ/L5HN73fsMG5mMk1nqCNUW5MHHMWDrJy4YOtUhYE6eBFju
eQ0b0/PCKXOsRuuDHsXCU2Nqs0UsqE8sD702zKa7XIvRfPjRxC16XPHIs0zSDAuw
94E8MfXaJp+0IjG+OufwsUFozhLpopcSeRRoFS5/EpG95FZLkNw5enat4/M4uGt0
LBT6D/EURrkTpWMJNzQNqOvUdJkG04AJywh3N2F3D9baRQy9DhYh6B+D7bdXABpP
ZHkcRqQNHOQ+0Ztnsi5Lm9q+QXB5bJaHju8+TjObfxUoyRU/iMl6kvk1FMIjvUBt
Sgiso4VkhMtybT18T3YOtgwGxI5fiCSsaNiTjDEXBTp1ux24MjdMyVjeRJi8NJ03
0QOGa05i4RfAEgv4MpgV3Deb6IISCrzCm5mcYNTJS26TUZliia/qu7wQU/Xjykhn
VXRpxUHSjf0mk+lVteLM1iMYIqJyaSasA8buyKy6SvGH5ZWaMP8gQi3JvOL5/Z8R
N1LkG4OPbAKZyf/q913Q6HmCtLp1N5RoNZIuxq6Ob0LPJ63dMqIG/tvxOrWp9zhc
RczaABDIdxDL0RY1KjJrl9Hk3Rkbyhd/X3Nw3ZT943kmo8kMOZHjjkYdcKIXEO4x
nwoszss0CFbLuMx/G9yk4nJ67/FW2amowrVAYI0avS8JZk6Qwz19OonbR4RNV+az
yZbjeXPES6kpk4QhpaLNOce0xRDZz39ECqQxOu/9HTaZ0Eya2N0E2qKVYQsFxjcI
d0QDgWEZBjmjXBqK3jqZaxCQ9muTZdd7paIVBsdVfV+2yydgvtmxaxnnpJrUDlf7
MhpMxtGqIx9dfpy7LdP3tfDMf82P4fMoDaoXaNa8GChLuho+mXru7mtpJc3+mS+E
KF7eZzy2BuvpDZv0ACGIvj+2fv97EfD8HO3+JprJVA6ymux313dQfG4ya+HFfBMi
e8vKahK4UCAy8T1mLwyKMyGupYKxwsaeLuXejzNxedrw+OUMhUT67y8q48w11Nci
WQHSz1YKTV3sVBfFIpcJFdJ1DXA1aSOravVoaa3aYAEIdkDZKMq98E3Q4xPVMO8q
EZa+YC6mFWKIUlSfR3xaTUB1jHFE8eNCcf4dgKPeq8BECXcf77lqI6q+ZpVwzqlG
SDuA18d4oY2/iXzakOP5Lv4+mG4wKua2BXWy3eLrZPPebs1aFFQ1X8f94kEKgPSK
RGTv59TFw65XzItHQQv76cewu0aRWP6pdzgVtdGssJ8C6UyzD/HFZHzVaTC1U7wb
lHNIPnfflX6eMm7sB03RJ6oMNMqIq+jcoydCUmfrSlHDwenimvE4RFxhDMx6T8u2
zuL0/brT5bOh64Zt8tjhcbSrUbILxJpJlxF88SxWvF3AVg1aYxzDEwCx++s/DojZ
PJzwH3DO/OJBm04q2TgyXUKQ3VKyMyGhxWOtfzbpNqIY4G6ptpIRpA0fM9OlMbCL
Thj6Ekx6JbEl8/5Kgb8XgG1HpbOurbTPsM9nzrlJWO49qRD/VeyXUT27pTfbxRzk
7suyOWvvXpXG1By23uof/LrhavwTmX3zPgd3LZX6JA6plJGZNCd5bDvF9sw338SY
iRzkjOGR3Ejjf3T/g9mnGDxudcA/SHxRJTEpF+Zo8j2XUXTcRJAHYSWE+qKuPqeV
qyvE9UXm2RhyWkEscyAuKYfGvfJZ8n0R3t+r9sBagZ8FJO9LThVeQ2G/QSdaafv9
vwMpOhITWYgZGMFK9A7i+n6qiCljLkX0pgvp9VZ7rXUInCwgm1IAjrt6AvR9vm9E
EnYjwecRwTwdw4St8Tjb4UZdKnbz4yMs8VreEBXUpBWutkMo0TAYVoIHP42viLi0
rSyElm551Ch9qPlX/tIyfC3Og6RpIyOaYGV6c5sKDKBkEYpMz5m8DYSHpDZZn/Fy
6vTZffxLcdAuo7YgHBR8Yb674e13eK47K7yYCa2tnM2tiOQd7Xw9aiPjpgwHZTk5
ZZQyTEtAF0htIEGNGR0BU5KpqFBraasCmv4pbWPm8RuCe/I0Q47Uox2PiwKzbXq/
a4chW07FG9E3+4++HHIZNHqMg0DnlEgYt2+l2UZy7vUJQio7Nqp3vlf6liE1cp87
sQwLT12Iz8EXrOBjQov5mHPufgAnF1mDBxlQeRwPNCRBHbREYQ8SCFYLrCLLjr3B
skY5osHfyOlczG4q3c1qttSCJuHAslwSW9Tt6e1T02erXRsRb4grXEvaE4SVpM5K
bYfs0rexWGfS4PErzAvBJEitz/VDPA4WQDhx5BrRn99MZKShUvaz3T3mdl/alFYP
pOsRcduCKit9u9NDmdKAMBC8InK3pipqIypsQUpqeFixrMR4B+7VYnp8Gbh9Os80
h+HnYvTycV8eMfVTFfheZdK7AYZ/7ngqeUXHU9ElH+DdQs0+O9m8G772wHTFpfEi
oIKLcUGxNlCmJq/rG1H9zzNp+jiNjFIjoACedqUZkDhDjK2qPRqoa0fjH5gyDNTf
xtQify7/nmmWHI7J/hTu7XsgnByEX6HvE5rwVZIBHEPmXnSxPMpvx2s0F490Nv+5
hZGK4SmcnkjauEVMh6F1gIfZLSmBa1aJV2h1Llrfu1xBMAkOHXbt/uih5VAk5oQY
agIIxSwSvjit/+z3zXpuLsyerT0GB01tbRvIfFsxtJsc0jMnzw8sI90+OltT2MF8
D0hHRzefG6nVQ7zEqArlvOSLlfx0cZZWGwOiBwEOcpQE5RY3CK+TytS0eUWZRpGU
poe3/HdqNx3/4fCfqpv0PtSLwIpJ3hqmCC/EzHvZBanDODHIAw++y3XkQaREv+ks
iS6lErseYL5vZ6r5yRKN9HLzBO5ot3tkbL06oIBJvEDUBD70zeThtDbSvc1/FqwP
6drUCuzS7fvcGo7QGm/SakMVJuW73NEYvA1qBQiLSkWxLqQraTVLQVz70hKaM/DQ
xNPeuZOyedSD4UGe/gP+EQnN8w9xn4glp0MuU152H8iOa+M4TI0UYeKWqM/xNPEX
iF55qXApykaADeRQgbWdPHJ8kuxL1oPA6jmVonCW6DwyJoBmpjAlhFpml3M9vEcW
T1NHfG7o6ZpMLGcPE8Uv2CkRcwdUh041UFQakfeJJl/+m8CDHSzg/Ptaf0xXQ6A2
V+Ggacu1b+UYHlBkSpGa+eCquZODc8RVTo/Af+kK7tgbYxLkpJgQw1VhbPstOz/R
dNLtgRa8HrxNXr1VAhyS8u7B0Sw1Q3903AanM+j2n/gnAyXsFU1GE11bSMB/L170
wVGvr8ItxPdvZ3gRJQLWU3TnidGgdio3i8qnZAVwnkxShPErX4j8LxGJo9Wg+iyt
O9Wk7PzPxuhilLu6jUnOZ8djMCGyv53koO0mSbTdhhzkpOllKhqoxhkgNegmzje8
dID4KKkYdR61mCH+OTLfzp+PbyntJvjNLLazrSDe+QeqXDbZYTVSwTJixMbeo52u
YENnczYwRHl0/ZwsxkTP18QiVEhQ4aqKB63MiCcOwfXfRg2vEPi5EVxbo31b5CY2
Ij7PBTSVusBNKZfO05j6otYXS/b0nHz6mdfvlzqfQ/i1KDZ+IvVQ2t6XspLYfozI
0YHSSZJ6zF7kb/MZ7SidS6QrB0/HOkwI813eNrtNcz8US6kK+xqfkJOQXIUVQaVz
szwaS9ofqi15RJJ7jjGonWQ109xKLI6Ip2BFOpeNb+2CNuur4WsVU9w+SV7q+WCu
NLTAMIKv4Hn0GScalhEyuOc+SpuiJ8K+l8Y88zoBAaZ1KTzK5nCBsuQov4B5tMWh
OGijhjn1clsH14xExGeEVDEhxQzQQ5QijKyU0QlARmZNgjrsArMY4zvf/LB8ZpHT
uOY+Gcz2RDhf5bh6XgX+WG8aboIUOEz9diqPZSXl6/f1XZl22nzMWEoeZldRNBGZ
N2RtsOVythiZdrOb56SzabyZBvqppvq8fwawZhvQbfdkzdrzDodrXcBuP1BNZC2D
r51hLAN0Dwtlk5aNrjQ8PQr0iWwsVIxXUKC0qs3wLvbDoOC24kyRaQgd2Es4JAGO
ON5u7KJJh53mm8CSabfTM+EvmR81uT7iP/FjlK2QPv6VE8P3SAhaUsFLyxl+P5FK
qUqOVQPxBOD6PpqLGccghnoGbRSaA5fA9po59xOikjYGEkK3XWcYDV98azNLbhVZ
+kxyyfv3BH2DKxXJxtqhbfqSztTz+Nf92ntD+8amc4TjH06loICh4towF9Re3j05
eCOATU4xXAFohLoE5RVZAyHfUguCcT+JGEZmLgJOctHukuCEPP3+0d1f+IihVvRn
NxmImO0FQK2ifOv3Okt/7kXpYpv2yH/8UYGKeGjpwGjtA77LqWUQwhLyWfvJTtCx
RSwxhHAUsm970SKTk7t/L4CiURmq33Eu0G7Bm/0ZKU6TeVrMLPyXN6pVwNeJWX1I
42VXa7BPEgxgbjzIf5lcpEGpnIqxT2yV+SGMFybkeO2Vi/3Y5/Rji6SVVHrTXmH3
PUrHsvn/Q69tBstP6VH3GZl3290oxM1qxI3SCODjXHQxHckBJgAQZ61Ml2822XFO
7p8OOjwc2PIIcs2nmte01p9jVFZFGiJAvg/ljc2M2pjS0z46ydWPCIl8j5HAZTH8
z4EJAMzLw8La7OY1fLDwalgRvaY3AAkWmUShakLuJP9D+WiOVbJ0dlqtDzckFP6E
mKaXoI0g8MHcBIv0iYrXxUYWZbhsP8q0iH3rK4qkzmrHfN7h3h/PTdkubMSAl/kt
PBfhrOgjmQ6Lgr+Dw2CLgGOToR2wV65grK9FKqbZZLNsoSy3NIpAhNTmovU69AHK
qYuQZ6WOOu7Lsi/oUz8u8/+mCiDAfhuxYF/UaAkah1P7aTcIYPBs86cbwkKpoKcg
zoCiQGWRBT1zMXItiLqzcMWGu0bps2Ycch99psEJuFmV8oYJOGlRSLGTXt7Z34lE
gy4CKHGkYiMNCnqEqEM8zj89t8wvaZfJ+HhhYYNwG5BxzRI0t0KGNgMk0RmcPxuv
gxDvnYPPcqxhgZrLFiqerO7gXfoGts8HOug86PKVfS0Cto6aDtQUhls30hZW6H24
wDbavrYIHZ5kK6kv1H/fJdrSgECvwVsqkPYlyLG/yrkcnVO5yxUBylSU+LPQbdPO
7fLlp0LzSAEOdzL5cx9STwrmS2FYMOQK2CWVQ/YCr0Rvx7NSiI6g2pHhroR810b/
NktKWrTLRc1mxCpb8IYtcwUyyWqVzV9eEWr7un5TmL7pmmo0LROBqUZsE5/Ns8oW
RATvaiuk95HnhLPQKKm5lJ8Pzihd5X7/zHWJ0EEb0Ttv2/nsrCyUZp8Dc304fRmR
iKtf1K1GE3IJeytiIL5Enh2eUm/BFaAimDiHRux+o97dpw/DDxfM6cBHqg1ziWCf
FXaP3u2ZtPu5NJsXzPwf4dA68ZzlxknsK6OJH+bUnw43HG93OFxNet0P0Z0IJXYH
oAk4+BGIsME4rLPNHxAMonRejk87DSRtghZVvSY991/pQSXdkgxAvK+dBAR4YmVt
TrDU/kwDOLjikOjn2ce0uGatc+hsi3HdhfAybDOY6xcBnO9KtEfR32btJz1X0ksT
y7VCTERGMufTB9UzBwWFbjLDqxa1CA3c183Rz/eTL07iJLkyt8dOKcSyVcE/WVbG
9d3a2hbBy6D4GVDOfgyc3kRvhGS6f3prGD21K7EjBTaykWCJu16QeUjNAaNHF6NN
2cexvY159ozxuknHP1BBzqENUoKDkCqVGzzEZDvbg0G4oYfyUfOdKCDDKKdPmA61
D35joQngWYJr68cdENLnFXLWgXXR1DHaHOUdTlkY4gVsVjTVjzFv9K50NC2Hagin
4/cNnB8wsUvx95AVvk09neohlLrxFXFsR5WjJwearKke27gmZ4x0gNI5s7TjBvuY
q+87rNeXy35fngNf8fLRuTVJ0XcFqyMEZBl/MNo1asgWN0ET5S8pA8Xc8jku7dIO
pScqXlTUETPnjJboUA/SosPZjtBbNRtpfLHk7kruEeQD9Ujzt0pB9BK6bwZJbSYf
7pXo+xCgkxTfyF+e0ucGv+wLT8LYXWLjLYf17TKdi6imh/x+y+GY9XyTyTV+3q7U
QCqXmoGi+G4IjFAaxa9zisLaxhXkI+fKl/wi2waGBBNvYKAWTGD7vKX1sdesG6MS
JdB+O+53IP0DDJ+1oLCaPbZy70vWEoNqhQ4XcweTBUEeeBK6q0mCy10hM6eh0iOB
5ZxFmXZpbIyH/uFT0z1Ds+C52IqpTg+VpRcP+Eccxg8SnUJLtiLnm94127E7FYIu
kuqL2RUNKR5N/TNT4kiF2vHnkOkJBhLA4NevGz7+cn+mREQFYP34dN3C6R27/7K/
gGpCUE27T0JcAu4bpyVVkl44yCHVJ1NlkgoVXnSPEh2vOmnnQf60Lf0Y1uKu8R5B
RZzUC4gZ/u8cBcS/DEAe3oy8UCZS1VwNa5o7H38QMAbTuOJNApC1gUvdePzIEX74
zs5QfbcDw8FuYjxxC7wma7qFsZpc2tzpoToNEkEb35FAv/3pnhDUwBB8AlJ4kmqR
BVMF6i5/Ol764jrfGeGOPl19FE8MK3TRxABqsaSEPFF4ndduUsZvD9ZfJ/G7AiKf
MdjZAJrV73b3mL8iyI+w5YD1vIo5SMrElwO6WuIkyQjAGff+r92kaRqadmKmOyKz
GMqFSkOKZdjtYwVrVWgXsPnroopln4pJcxQSWIkzkdxWAyrJrU18RRPYL0nMrI81
LN/B+/l1+SuCdfEuzaoA7uA41MVKOwUP0ud+JQ6fm79ySCHyb9hYpCtD3j7K0J5m
xq6QHJGLHquqTc8YxrYhOVWKhAM/ooZ9N8eD1ZoC3Usmd7iSDVVhX9YoDn+AdSo6
N0JL6LBGl9w+Mqz4SJ9nx/VTse8RAtyqTkskfXmmnxIK501IqwTgPx25rGTcgoSd
XQ5dZQ2TBz3h+WuMUyzoSQNCvu8zwVAToyuwWcC/uLiS2b0Jz+5UShi7fzDbx4IZ
JpkLtekiGo3pnsAfq7vDXPtYgo1dBVXJoGx9lITLQ6xiPNLnDjwsqmStK0U32Ydr
e+CnSwyD3j6hEIxw4ZPmnkQtKP+TnFv2AWOA79QCXzU1WreP/N84A4CqEdosuE1r
/FXSWDaTFgaPnXGoqNVmiGip9PJayIHEP5fJAubDbreZUWUPsEP74hKNvcn9X7Sq
bhz0VeMixrJAIpxWBPBZpO1TvDlZ58SwLxD+8GVt/RzZAw3Mybk3WDhNBRu0BkIp
FkfGSnGV2ys9vyQ1b5C7bdcs/WNirq9Q4jxD11nlp18a2iU0Cm3G5HszXMwvMaCv
SWFuwe9uS1NrjR5Fk3a0TNFZPyyqvh7s1wjkz7ryb2Fn5jdmEjclyPca31ogLMm5
TdlsPf4UbIqwqpiRv0BXqeDtIz+LsgdKbKBkes8EAs1D99bH2wIv1SHVvYAFhDc2
LAHIerWEfxNnPbDScVq6lZ4grEFByf9eVAc9l0QxM7hz0Dk2vi1Q9rQ21PwQFAjp
Y1Bd2Y0xOKqc63fatIYhBgJuG+e1dT7yqt4Wz8Sip2Y7t9UO7M4CI6vDZPsnFH9F
H4UDaRsiTDyGRgZH0WpH4W7OgXVLWIrfqZyF1kPJIlOVqCESWPigyo+lQzkrd4p0
xyyopglpmXPlMZpQef5f0pbwVOcQldy39HpzBu8nKGCdGOf9Cr3ToiRGtp2kX7Ue
Hz94CpL2cTlkTeQpg+GHE+oMnyS4G3fufuDyo3eKbsDZhM1yaJ+/k4aHQVTX4lKZ
3JhIbnBoUlD5ShM5RrrPsJenLqVsCY8JlyjSuPNa/phnFgOYVw2iiSUEUfeDfvMV
9bEIesRHGeoetJrdTMD2U53woAMChTeajLUcgdTfbr/8hLSHUVd7tiT5kDfCSqvM
5U4jDk9z9eorFrpPp3YG/dkikk66eFCXvm1aLJiu1ejvwk/Wwwom8uOGEhBQ75bq
txRe5pRPqtk3ItOZWjwcnzQLqAcnnuV6L+cfBbHX9QI3LscJPrsOwqlDpKyLJ2L8
mkOvT7jayvWxfuaKtBtDcIj1BZzthiqtdql78Pf082+lVwRWMOLTPa8Hf2dPb8cw
WOOLljEGwiv5a+WMOYAc+FMEVoDItkAKZIXmjnEV05bt7EFc1Gdog0CTTlBJMhtL
kPWrvWntlcqycFDM/N1K887pZxbowW4Xt/meOHoyE8hrJtf7WHp54nNzpjDWFC13
CyKTPPzSXMeLcW/xW7mSNzvFpAsoODvAR7MfW12T31eAeXv4WfDBzT+YF1vg3FGR
KOQ/M/z6zf3ffadmAyF12WBNJqih8H6DcZFB7LLJ7bMbKgRmXNbhE9Y2r7GeWFek
Hdon48nIOGut3oTJDT2FjOlFLqWzqlsLUOWiZwEDWCnv1wPrP9M9gul+1dUtgDNR
mOUgGMUtzlt0a+aUCoA6Z4CZvP2tCEAyVE6nZoRkZ0FgDKA6raqhn791DD8viCm8
18j7CqDWk1Ux1JSpV3tLP+WvXo4iH2eyXueA4OhLVjL9516JdUfQHVlzzhTVdKxm
X/6cVScb7t5kQeaSTTrPCIVkrqCkNwAaDOOwfk9+vPBrkTzhofPWQN/QG3rd93J3
n9w0+qIuxBYcFeATNLsoMMLGtvzlX2wFepI//rvEh34wlsqQU0Pc8X9+VVpEJF+N
U05eOmlNPOupGfoCfhC9Apl1lyDHFow5irhhAh4pwCpKb9U/CCFzQJjlaNHeB5Sq
nuolZN28B04a+uBgyDXgiSNDA/770RiAx3zQf4CkvprntdWAOjh2QXSgG8Pm3dM6
9hGz82xmXSsFBnN3LkBhWnrOs5iveYWCtLFsTEipxNpEtL4AB/SHLL6u17d8jkzk
BIdIjJF2jfdv+JN5BRbXm0gvkqBDH7VXTDLtWSXIzF5CDkY0//IU7d98AN6MdqMZ
UFkeIK4pEP/SfDlI7WzU18LYgZj+CS8qYe7S/q3icaT4p+G2pXC7QiJOcr4U66v5
CEjYv9hGjF1Z6SwKa9d3zB+J2vRP+e4Zi7GPAVnEd/J/0aUSUcSrtSmg4k+zN20w
+7bnuU+EYLbf7L83my5g6iPxenr9jaXyKoyTEobTQufkqonfOIPF7ZZXzfRxNxME
9EBGMk64/UJYaqTY4AM6iKO8usnejekX9p00FJ6HYYJ3oPTwSMVQIvzGGu3w5sPg
204Nkvqn20WQma33Le6/uifkbv4bd9L1hgxZzdP4+rp7zcy7w2K/tI52eCXAKrl/
ELnz5ysDI0Bw20Ga0E3y9NHwBpZjjVvqKCBiUEaf+CFQTa2rEBVS+hr6V//kj0w8
9p77WPkUHRNXQW/WT3Z7fDuStHig7ndhx50ue72B3gikQxBLFVWbDIFs/A9YS5Ao
5pElMNPRIBO0KxL3f7P4wg1EhhFL8DeWru0d67nYWU+DiEM+ueUOzSU4ayMWcg/r
qCBPe9gAmmx7cQB5x5O5vox7GX93KvylfzIBtAe/QVqX5hnFca8ZXI+me/t7ZRnN
LkzjVAYIAEXUSkYCpWqLmJfTi0Yev9s685f6J9nT+pLNzOwaa0W7hHf+uWpiaSf2
0cbUjmc4zt+jKtBcCqUQpo/uq7+GpmpfnikiFTKdU22IDAbknmvId9llyWFKNHNf
WTIO7Y+QjrhiRCOAZod79YV8fQkMVgXE+2e5zDNoe5CmXJiMuDMKoV4GmRZ3cg9w
dc1xjeHd2SojdulGTkeWS34t4xAdf8O1Uq0ZwMo+E19Ilz7W0zKEXu8Pf2sFPJgS
S03cN2t1WS6O8BtqdpOC5kiym5FYe3oYPuAb5k2h8LrtoL8SrhlL84Esbzah0p07
ROVbPge9mhrVKYY/nmRhGNG+xLfJPIn8KKdzj5bUozJdMvHHOY/0gs/CJ1kwYrCV
dllr6ikrDny49zQNxZi+n8mYnYEL5523zpf66oSX9OrmcOuSBIlvPDVteBcD/76F
eOVFhc2WdD6rc3JYnu2I0SyWxKeAXdSOeAV5fbCztUZjNAGOOmzchg4PrdwNLFF8
RROlO4/iie4Tzd0k2BGlk6iKj5X4tTt23c216dz12tpXRptmi+jf6CdV2YnihEAP
WroM6O9vtbLyVXuyUE7VpGMtwLlaLzwhmbSAXvicdV5u9Tekd5h81ygCAIraZDsG
ID9NaobNqFJFOir8xgXnWYiu2rCRb9HREDMegjwHDrNJFiamtx4PbdnaviGYURth
rarAMUS5mDxL6K0HByWd3fj+6qPGPX7mWguew0bxGoSoW7IsRASKbE0sLID1jPxp
ctsHe9cDbgacMWLThUeERAM+KsL9di/DCTGhx8n1xruiGIewtojlR4jdAn/N2TA8
oZ20Hm0ofctOg+JR/iS3kaj53YvT29qWBzvF3+AxP0zHlfUz7q35EcTPxOA6w3n7
vI4sQnO9vGZTK7TclRYA1xYVdSIj5DTR51dI0F8eIGAIDghlHNuZqlpDCWwk7O1o
1uJeswc5Xog1Lpt3wobojTNnfwqk2xnSXDicHST4VQDFmmQL3+uUZzigBsIA/6KJ
TEls7dg+g8ydZXfboLuhKp/OMMbnFVFYb6iWnu/ihmd27f7d+YVytyjglg7A/p51
0Px6ebVxipEKmQZDnTLLpYq8+WFGWho5RoKhYp4OvPGqcb9izbzbfufo45cvwo4W
yQM4a3z2DuNPEOgtSdiOBgZQsjrNJROVBv6bnMZmY6j/NsPSAum0NEYv8aU20WlS
78gZcVhQYYBMOR4+4jgHzdtYiT9JafBYxRonQxFS3d+fZyvjts3THGV24bAVtF6p
iMhxBMYBN+eJy5LtKmy31BpFag7e+TDfcGroZmIgkyV3lrJAMBvYjJQqsJuifat7
Qa4Z3tHEuBg35DLrjQLHtV2YgKL3O29NWcX7s3VCeXzKOpc0px/0lbmo1XJrRbGe
KmDttDA3EilmMDAHxnyDiuEKtL05EDqpal2lY2p35gNJgLdonDGeJtIgtTm9sx6y
4lhBgaB+UYHecwYzpUxgY6+f+0R9vdbn7d+6x/Xf8rp/fqnCiGhKXS7hjO+gaOOn
K08SNcZ7qAG9yHhzjtoEMXWENq9idcd3yBjO+feQhX3dZfr6TQtlzgPOMpHmjamp
6dEG4qfM8aWCKf0RzjsQ2kiw8gpNpaw3G5jY0mqsu4Nf14Sv595v/kqLQi91rQhB
/QRS0LGxi9PFJDDypy+crWSPTBjS+74kOxTlwpAWSiaQObxudJC+B7PLms2F0yPp
0ufNrXW/QyklfNVy8EA4lky3uO0WLkdyVYNHXXgq4ILMixUASdAjEqsCYsWzWp2l
o4jMvmdkYlp1HeygjZUWjwLmLpkyRbTin0t/5cWzz+KypNvuO7vsINpyGWfKe7VM
1kDDt5VeOD2lZyUENOCw1h+hyaN0VDpIe3jqau9zKg3RP2w3jVG+S5DCvI98l9Gu
COgYkt8gK5Kxx4bvb8HDhpeuuH0008rAwVjuB1C6FOgEjPEZq+E9JtjE0CQLAIAn
SrD9eXLvTtgOji8uFCWvYhmGQbe34oNjqvsTuYE3EZxYiX5+6DOREJ5vu0XllG04
NaPUehrvslmjsQ+RUvsn1UsKrFl7rE0SUOC2oJvSVPrmty9VZ5Y34cbl89kpn4Bm
Dx4I7Xjvec0ipQMwHnt9+P0HeUTt1f+NlILuCu9DqPevi2RB3h+QSN72uUMpDSks
4LwOz+CmLp/R6nOIvTCZqmpraJ3m+t3Ja7cZ0u58GyxDonLLGOS/uKb36wJ+xiuj
VKDbMHYp9wvUC1rNccAkrAMS8UkC8MQ1Wv3JXF4KgwCVdY7H9Xvx2nnxHuGfjIzs
Fz4YPWaSTdnkUk3Qv17wF3HoGKWmQc4efGUbP7ozxv+XMf+/3h87IXhAcCoji+Mo
VKvcORf0s1JuhZe/kBTCCPfh25475hBLsiki7MdWBWzZtz/0ezSkIHp1xcpuADt8
DTzilGp/NN8TBMImoiNYLX9l6DnGSOU2xGLJ2sgcgtGYA2A8i62Y9SnC4yDZ8Atf
bZGSoHhCZkrNFL8FcvTHj3Q14bn4KX0Bl4y759BAaiptH5l07mLURLSZnxJ/7dFN
FJpRAI/nzBRqBBY/Pbpe1OW4zkh4kkX5CPqpPmZUTMbFoePnHMt5fANYKn85blxj
jGXL0fDwvqBMKSXe78Qso5po95FR5jx/3FT8dGu4wKnQzQvRMXFLQzvnNNqVIKj7
Z646PAABWNqoH6OxRB//79lBrHk9igpYT/KZZFaO/4LdEnd8m8B+zeCHYRgPyfr9
75sRHzT49e0AfE0RQyheksoeDyYQ9lClpWMQfmbzolNil7ComNA2VnrsM1NHLuij
pYNVtivFreEKhf53ZuIYFr339uZjU0AygKJ0B4d4BJcFBlwn+cPdEiBfXxQ9miJM
ZaP7hKLFx8Hp7QRfFYLkcfCbp6/BlAA8bcWlpGw/ptD2dqle2a4ciyRL0F4zMfzT
gbjDXz9RCBsYtbEbfmY9+Vr6kRIMNdlUUyO+rPjr7r4amtPM6dNHYftr/rn/FZoi
CAUtx0Jrf8XmcWPkO3eRJ/yeazCbR3LNOxwPM84efnItFDsC0ZmtgiHckJpMxWWu
QzuhPO4r9UBE4NhrlCAFflLT/T/OqWYGHqDQIltZxbHYoAxe1vjQ4uyYTRjUcJWf
XNgjSSaU1VS0dXcm+5UZQz2F3S/rd5mXoKNUd5fC//aHcngoGgx0WaiHJQvpfxhA
TikXJmYDzxxB0BrFWfLnsIqt0Gg7GvP5+TeH+mn5n+p9Issx9APW1kauoTcNaSyI
9yIaWHq2tdtsvEUQ4yKIeESb7+4jV0TU1m1OFTh6uURcHio5vpHAn0+Pw4uYB0o3
d2M3pbJZrdH84NXa6wfYwPrheClulleRNWdupZHKQG16CNXQf8DKfDyUbMiamTbS
SnmSYXDODZrX4zp+5n4bJl093b9r9eCybHlO/JF1qGW4X9s2Z0nYIEfCPbWzfdO6
vlnp0O9hJatUEDaa131K/Z+jtrkgFiBQC00yr/o5XP6r8hB3NQxBfaPjQebBO7aI
dRYZmG5BUnbMqRBBNCKlOfhbEFHuU1kr6NL8jjM5w6WdjTS9UxPi9OURFVkkktAX
EdvmvxcFxN4zTvBYD1poKnAbbfbz1HchrUS92CTjYfZ02meXrMgJqRky92ERsBM2
D5Ou99+MNu6m0gwkKpWjYgysOR/vt4MkUj2EDMy6+us4dFc92M1rS4+gSDRN1OGC
3/uS8ZVsQf0sMHstf7SNjfTYhOM1L0PpoO7/xkwzvXth/4wNHL7RjKG4tuu3QiGT
dH6fnVV8nM0wDikBKtoEygkrgRWnP7C0QLr29s0WAudtM/kiASf5IvK4TjaxBKJe
VEZ6wgqa9rZzu2DsDd2B7arLhY4dZqsOzLUQzqnHAf8K+6efsNaksj4m8VCzdywO
aMK8neziuqIneohpxAP1aV20AHMFN/EkqyUhJNWHYqi5qv+8M9f1cWwA9T+dTNIf
r0+6mwov1UVQ1P0KAE1HxcPVATshXn4QvnL+5QCZqzCWRlkFa0zMTx3+fqe+Iqp6
8r6tFQo9L/INOhVuxkNzWvRXLFFCbMEcxDJPsAt1Swq+1txkjiEUwV3SOoactHCg
Kb8UEByULbt7t4fIM3WgUYr6BBwR5JynqQZkFq3raoWGyTdxs/WyP7cjeumWxiMR
vrnJg91gHBNLOEz8a0WlnSebBw8Ea5CfWHc2BKF2WWSHWJPmNnQAsexTg52MZewq
tb/GaB2maFjIwG8iG7BoKPukJLiEHrioA8jDknWR4tVEfhI81puc7UGfkonobDPe
wNZA7Vbi6BaZd2YWHVQOt0YrsAVO2ZAG45SmbPvonrhmm5hgRr677kz7O9XlPvyY
oS1thu33k26BeaOWANSJxBE7WDOVFvLCkYu9p7yV3optRTJPYK470XUuk+45wXBs
oV+HNxZLHVLK8ZS8ad58Lp0vXMFStUbbg3exQVHvOoGtfymaqdpr2w1OnQhKKrK+
9oYjL7lbBsqdfZhje6RoCk142DiI05O+519J+11IGdT5lnpXauSod/4IrTMi1e4l
BogY2xPOmo43mdQNy/st4XUbACWYvZSc7lsrGmxhjj3O34vajpRb9cYfYAUMCQQn
TH1TqZwMwJJtqAZfOggGO/SjCNNP1oQ1My/EuiaALfMe8/kaJrVQlsMzHt+1/l8k
IrKWOFssO1z4lmQg7McyEKKx04KNW/tWCUfk1rmdLgU5YWEyqjEbdUbq8nla5qUE
yOshbffbq097xZ7QCRCf6N6d2Ojr4E7QeLQJV9S5dmL/EptpthKaa0H1lkTkbc/u
0mLHK3Bo4j50A6IJR9QXA7ObYprUEciLe80SXpsSewWRgSFpxbOPX88y5vUAqKu1
TG15EPBVel/ZLQO2Y1DT7SZkrFIyYogUA29w9iYfW7OsjOgnHt3sHQkuqyFM/rXu
O5IhO1wUHXwTJjO/ZaBHr8SsAp2ZmiySD/KvVl6uMMxxHWg04FuHJ/YSup8gGYFd
2gUIJjfVtJC3JhFMLlYS3qd8DPhkZ/AJBro6yFWoAej5LA7jgKS6wUUoaOLXVNth
2H/yW3mICquDR5oQRvpH5Ae3R5NJXYwinU0CICyA1P1YqKOXHVxclM0LX5X3r4oI
bx+wFkxCEWc9TFF9NOyxLhpXkjAfAX86iqdcQU7O/7W/fHO1uJ2meFYys1BDvTjC
YjEURHx0R8ahFSIWf1Rav2heAwDFrMdXkR6XsYFzNIyltlLnzXTBehXznCRFiXNg
iB8dA0lczqw70oDaWhuKS94g/6aURl12trKh+bm3UoFKhMn4RuYiHSMhdqtZtuh2
U9Uj5nZIKViv7Ucjj0tXkMYa+Ylzz96bV786cBPusR0PGvocJ4wg+RzArj4lh/5B
opZkiy78LGr2rMnfyHx3CqyoofZZzxhDJdDsvsjSNGb9pnuZAn023SO4Cv5UJ5w/
vNmFqQ0YS8Q7Q3W6Q4kOVGn1bjYGToX/F0TbyK7z/BRQZI8OODCCHvcuim6slPpx
ExyKAncWmbWlt8qdnrHUjKQUxMpBbMQ09svumeGlQEWsOoryu3W+J8btQBQz4yij
aCMoeoJdlEBn2FVXPZP2i4+IjOmmdn+rMqgKbAofvRyd56n8jIuofo7m7ig3iPuv
mUwFPc0id45lThnMYfeYPr4D+dKdakWhfRmTOkwzGkbdvn3KO/JSocIOwQrUHyFI
b16bDUH2K48zrLH37mCNsNKbl4YyLdkogHqJxLt4kjk3X58DIgvVYxVyphstYIny
YEMz36LYY6Nhf2xAtgBNMoTf1moDOYxYBk6cajwlqTazRB5tws68KvMwn0c2J0hw
fLUdFZbzCLQMog3Uu5ywPG42gl0bujAqdCMjNfpG9EDPQ8XCFU7hfZIoH/zdZ4GW
C1dBpXZExcsn0K2tgLm7ljlkzeU3zr9UQqm9ZP2bKXRJWJVemH62Fkd3TfJyDMSn
x6gbT4znc3sK2jdBVSUAhN27O30l92eeHfcytGpaoOh2vsvPrytQ6rtXbm680aJH
e+rS9IoKuTOi2mPW4RPwZ+enfLl58XOZu5gm5+P/q5NSJjwMS0HW3nZp3nhI+M8u
G0V3BxruL5zIs/PqfSZumxJVGl5aryX9mTbKrxCfIMPS0Pli1k7HOLIH7k0ZTw9k
yJW0rQvFzCgHTfzBJ9bNjGfNNtQYkWH01mw1CsQ93daFgklayFfxlDuvKYdaVKKo
fhHd3D5WyaUQhiR8vUoazuMBcekurlP+BvsaPFBb90OPhrUkekZn+N7S80VneGe8
FczSaZt6Z9W13/UUrDiqVacdZGCV6XpqikWXH5tYUkS+aWwF5z7/pL3FKg475uPn
pVM12WJT6PfT3NjLJYi3sqKYc5FZcgTWpD3hP3Di030bWYV33dVybGqSusx/cBfj
LHUaahPSgk9l9yV46z/KpppmDeicLtoh+7+IiAyAB/GG5eZ2lRj9f+tsttpHeZPR
q6Rfd9uwViZZ1nJH9uRnnuTTo63+dmGyaiy4kxzMPFUlq0n09vrAp2kZ8DN9Np5o
fc+WNG9cVi65UzBIqVQFdr+aDrY/DhQyd0hYaPnxaGRwDWkXAeCgUF77iYZxTw/n
o5FaNTLIrlFc7ObD+CVY/qiVJf9EsEL/B9zi+OoL2pvCeP9G2WJm2R6ZhMqO3bSK
0pDEBm77B5gHlEYo2uvGdtU4IINPDHKpjIidRc0xYBjUTEV5grexrx3A3df6a9ty
I02KuPWMoOc72wVir8EdkwxBzYhWuL6d7lgtebUC59iz8bOouCpmhNfhyuYXbBo+
ZR9OlzldSS4viRXIq0WaPSnOzZ58HcicQrbFdDRkcRufyKCYl/xqKbahoGBpgBA0
3jCsWNZuWsf4yIPRmiNQdEHjPIf/WET3fot3TRkaPE76B6KDJxSSelO5fP35PBI3
bYHWRVzKaR24jqa9n0BJYrWH0dZv9sEddQkFOEkJfPVKeC6gbkq7coUYBqRXQI4k
QHExN7Jb1WS3znJEIecYQ5IUM/IVJU7WDqEIRNGtCzUmBLBEW4YAcSNTSQLIgiBA
A7Kt5jCRVBqfJhvIYB1PqNdYf3/HcxrH46CmvNzQhdQGgVnZZ/DTDxLZYrtQtNM8
9HmpJcm8bEeXNoUvux0BVq7iFv8c8H8R4avZgQU7h+MIAKeZJu03S+wGZ+p7BDI/
pYHgeRt7O2xyQ5UE9/65WVvABOll/qjHqG/t17sT/pX8ZhZGd/gTYJsUtk6M9YLr
Zii3evjSEdgwqSiOx4Kjp2T9ux4Q10gH/rGsC8ycifnLpBMyd1ed1VQhAC28j8rz
E+qADtkzBomJFrKEfsWPEkh3U9PJuRs4XGU+OC0YgkUCW+cYfJoXa1z98d0lCQWa
WIBCBbU2UVfNhLY8TFi/ZUQkYm5pwhpP9q4UHwET6v8+hle7y4tuCsmeJNufQXs6
okENHLp1i1LghyB7bMLfSDgylg8dAitLpqe1WbLLSVpK9frkrlv11TF52UA82t0x
j2mQNxzBKMy+gIuCPy3AhHhiB/BnrzF54GvrJaV314TYtTUsES69I1sYsAWl0Axq
lw3d/GXTLnDPsl0MM5M2GeSaEbpoJ3Cc/L07ycXHFAn417m+Rp5SQjLwiQZ8S7NK
D58d0WvsID9qXPRHvz7ntkSx5++Aq24tBcyJ3foejH9Dd1x5/GpGFT/UasOxZeaE
nds6WtWLj8S0f8morQQkhchLjbp0I+rTE76KcyW7hM3kNbgK8KTh02FOTEVVyh2J
bvFaDHkdIE/jk4atPqbJ0bMh8maa0BSt7Dib23Fa//lIIMS4NsT6CgdsAyeQK9a6
/W2Ps9d85sdQwAimtnVZuvIfAhtFOVV5zTPFsmsAczGb8cO5YkSwTXEcRrJhZGtZ
Ow8RtivrWVq7RXD3+1HZd0fFbXPbg3q4p6a1HQ33VSY1WuoOlvP2KGvG+V8ht1GY
/9AjbQ5ixzEcpDFTeecGTN5uvbbPhCknHW3mRH8fy7oGqmQUOJ5Qph/IYwAwfuF5
HxgRgTgPYzSYrC7Qw9m/bfUln+hdU94tYK/Uxs4/P3ewmXClupZ1KAqMrph7cY53
6i6YFv8zwcsYlzfBPi1YuzDmgySHRgCJTlulCGniisXA8CVdMSNCU7J9e1/+HP9Y
a/5+sAFe9hedVA2MDgHjGsj8OiUCOIhpM0y9Dtoq8zivc0wPlA2ARbOZ3eXVUT3A
jeWjxYjkyYVSEZRY0xJCq4uvbsNL7gVF3bM7obUrSxspXqOvAKhwNSlDRqiRiNIs
Rc8kxuwRdVGZeVgN6ICDp6GC7RcI3quXdbdJKO+ZpqBAA7CZ9hxrfj3Jp4Fv+99b
VLTaDV/owuV22wEPZnCF8Vc+7phNNJJXuUiZbcxlYPcgrqGWbLEXgjR08DzLmAMY
bt2p4tqaByq9U47j0/yTOe/1dR0hOjfEuIAF6pH/kDUmjhHJCPeQQzxC/0d7Xpfe
HH+HBTZG3RP7e+5H9AvIlbQk2lph+upaCsHUkU4z3i/Q+upz3J83gEXhpjJG6lLo
i/lASY0K+xOo4uOuSEmCJ/vIHRqyYfsTVcU3nbwsxxGgmaC4aGfBDxXNyg1iTpyf
LC8uJfy3uzvsCih5dM5eFRKPDEEIahNq37Zr3hiuVh1asn+agWQrePoiCJeX4dxU
p9ZJgcohxEIGE2amcnknh3tMVAwtu2JfgznVgsKB2QvAcJ6excGizRKee9KG/GjS
bq2oSj9A7fwQeaZ6xwmjlVlLywp3Gkavi+3/I0Z71RCwz6bY3dpwhtNhS/zdpExl
zcZc8mj4TbPxjqBC+y10p/mJ8Z7GX2bMgcsYuLfccUTzW3ew23hrI2O+QNB2QPJe
wCWp580LM6vlqZ/SCivqShFSxzvg/b6mggfrSlgWTA2q0VvOwePog65lwGgDEvT8
rJKbNC34qhc+lfMUTFT8CKuxSPuW36iqnllDEQv+a6fwpBpcQtKkybqX2JzjG13S
F8vOUOJWvHSWuoEBXteu6Wmj1WP1UrEz0cKdxO/VL5i8k9G7r62xRab/FgfqgUYP
pdmqV7PyvIVNq0yTWPzFDY9IIimE3LjbFxqCKinizXmhqBdCaw/W+XHnrNcStFj7
nq5J0BfyJfaLMCK8olvMGT02lxLWE8hl6z4NkDX264UUM74VHb2oK6NXQAymd/qS
Jt1k5aaRvyka/JQ9j4Ev5yknSe1R2cLq5Fb1elclzdr5XcLyWBaIIfzd1PytxrrC
xV/TRI21JrMt+dqHUAdKz5WJO0dko/TJi70FCLK9hkLxufdJjH70ogvk6/YmTIoP
pd9GKmxl65WUk0bHMfqwSj6Bpg0NdVVTR9pW2nKThhPgbCP5Y/islUSRrmAFLcQr
9SwX53kl3DcHFpl1L3I+cEvpCRjGWlPt/DpPFAppBLFH4gqY43DgPRMNsu7eNJHm
T/Mi66UoNkRAm8lEpTIz8wFbVGEhNW8oGQQgKSyFGzo59SvDMYKIheNTY3BqvvHs
zVTWM834iWO3gM0Vxl9C55bxgAc3QRKpSt8VuV3qiwn5/EkIeucuu69JCNJhyuau
FtXHQBCXRgoTeNSa2lLTEEAzxHhWqoOtU6ofZaLFXFl5a3COA5pTAbnWwQJcgA8i
x10803L1Wjo5cNJcGJcYXs9yEqNMDLlwOA9qVlV8C9Ys06c1wpVTka7bf1TXn0GD
eUm03eKGBkWxuRLkDIQMSaDd/AcfvqeoGwYEvnEf235Ox8fjcowFd53N5bvQWCfY
RedQeehnN/Lwt3/+EchufJwtnFt0kY6Ptq6QcA9FZRabfsl4ZeI7BKfSryvULfdE
jOD0ZESbOPgvwPPRDpxpNc0U3q/k2zCgsISQhyBKKXMFnRhRYf4ys5NsGnWRLvrT
A1OCUx2xsN2yu1XUCB7TCX51TecuhjAEGeNdZjgpfgxVp4fCh8LGKKVnKuaVhigc
o9Kssjfxx+bwp4GXl/gT5B1eJ/0FtkpuuBgSOWm1cCIpUBjfqeZ4oe7yAV8jhSNs
ZDbJRzNTJ1XzwPj7FSb+m2yD61Umt+vaZWiWw1LCJLjfw/zVpIrWPprzA6/vzSWu
IAFVTooO7sPJfYuS6npslyGAoYPiC+ueYzi/hY6dwpN+GkCMHZFBELjBlaGvZpda
BHXru9MvMvQDHr0wHewGlRoFcbM0xVjATMubCc/QuC3Rct1sY7MpXf49H8jblGO8
m4hkG/Cod97BFrSoCH02F44gmCiLTkONaQYLpNtT819ibXl9XQR7ti1X+XIfjFbl
ENHQ5uzmvbR92tzhVIL33suJitPaB8L41b4l8VTWkbo9Ap0JmtG2OlyRewraUMCL
RFfsCyg5HxSwxnG1jgyxvrhDMgX5WzitUlSMdct3P69ksggnKWLmZYA/trX7iNgZ
yvPF9SkL4u4hnFDC+zw36HJoltxmR/G/ph7gs6tJkba+pFmDudrzuKqhhQgpbMnZ
d1FCXqcYJtz/mMuHcEMH9Bl41VW3H6EviCGr/E43HD9Y6fYE5l4a7sEh+NcANefZ
xoJtXchCQH7+VyfDoOlQ176dwZIRVv2zxOaNmCK5DuVInqENUcKsjsakrPxUsIal
IrIQsRqTyJk56R4REtjWidfBjuwFJxRddbsVZvFVFdUY9nS4WjJJdy57CUXVnr6V
ncc7e7ZAALloeSv9pjVPEk6xRGY3hAXfB3O1v6oV3uTrtUZdiI6T9ZTQuZpbejkr
E+EDe6lZ7Zw4+hXo9U8sXAeg5iw2KzTvcokilQl32Qy4F9+n/OqX9ovgfYt8atJP
2f9RcaY6BR08iluiR//Jy/yva41JqUfULhvnnb6LGfIWhf6oGi+ecZayFY8gbiMY
PQWXCTtIo5xakhAYHZSPUocp4/3QSZNdSIbzcaCjJYkQk+lAXlnL8a0fphfwN6/F
wZF4k28/d8TEUnEc33d+Oq/UnUO+D/q9vL6VKAfZgX1M2FcaYeGR1gqZDHmMs2Qi
7aulrJo1oxSb7CvA0ff6XHOlwj+KfrYdLwb7ZextFxYkxOPHlvU7JnwBeIQI1H+K
aAEPHhHWaUcgoKjR+BvX4t+8aa+eItkKHK3TJZH4ux8EtpUx7yHjSPtZx1bsw4iQ
GUMai+0fupCPg0EnwIO+zioOgtZQzW66ORQHyNNZhmldqdBF884rZVTvUumGDK6Y
SfDw56SoxmTcOz4IgrQaqgbnBQxAABMpTlwbxNFPFfcC5cvp9jYPDss4aGg9b5Zw
hRSE6ryHHctSxZxwKzQSDOFveFZatwt+8IuRhNjqzkYaOW+fKSnDKM/h6nO6Sa7T
tgIQ4DWMS5UuLb/dqEHoyY2FdlIiVxBgKIZfZuzvJGnStC378pV5f8a6/Jip9zTr
ZPlDyqNSwSGM/a4Fx75PWckxDIGMao/h7Bxi1uQTVABNm34YKe5Qz2CfSiYf+BKN
xNDUIeXhgtFHs4Pez6De99vDzYj9XMoP88vgTpyRYJoAN1kCFMzc+EhkBrDbsaou
j0xgBAqb5SynKOzYnkhluRgXecZWu6CPu9tyiz2MRcjjB25hy8fH3uE7JM8VSIMz
7IqptxD0M9glN51/wzYhzYmaTwUK4wbl4jPm+2gF3vEoZW6M3wyudWXsEut0SAaZ
qn2ICpxIJqFQqNpBOCAbUQeIJjhuIqjnu7l7cqy2XELAFVifeXRG0DLhcrhttXDQ
e5efNGb2qFxO4gH1UeVdEGHwIIVca9H0eL4eejmuyMJS0eh6BEKOTCTSIDJ9mEKX
Xh1kt3b4Z56phVPIm5iEmGJDICtdHlpVPy1FZPThvT2KEPDF6NfBGESiwwyQvthv
uU9xWY+sSIYszuzP/+Qd79wDHIWQ5u9MUInaY7VWPJi656tO663XEuz7jZj8bAZv
Zd/zcv1zlG9YHF6uPiXxDHm3guemYEnsUIXAtEZkYHvxm/vgqBDxZwph8gVaYk7a
WJIhTRy4HbPljnNeyv5VoSwy7wLrbgD4rqzva5QxRxt9b2ESfOYLUIjcYIpzr4uI
NqvozCATIgCIuRcMegtwTuTQlJRrf6SXVlHxOeE3N48qIP3It12R1/3VtSHofRVT
GGQCe4TydFXYMJ7oiyuDjCY9CgSiJq9IC7j7aPg5Ar4gK69iPOsA1Laj1J6JzxEu
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OwhNDmwLIljDSkXkzPplNSub+m8vAJbNFWNINF03m5pJ+qwlrs/jJHLtUsto0EHq
IWh1ECFu/XPpF5wqAc5MTOEWR/YXNfrONOZcqRv7lUJJChMTZSHkxCoLpA+5gM2g
oaoRtfdMEERACXRlr914QAy421php+MKCuQjz/ksCHDOlGscOdtl12/GdEWOfGXd
gi11W+lPCRaOIB/kkYN40cabtoIiFjazjPJX+uQYLNsr446Q6ntvRIMhE/xExhPu
JwTD3RFdE14EtNtUrXzHw6Swh72/Oet9r08ntibb7Cfm7Oqjt84ppnkv2xOMeP2j
s0p4/UNkiddnL0XjvbAQkg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6800 )
`pragma protect data_block
mjAqpDzK9PFWeiN+UuYHE2RegMCFHXHSoJirt9ySC+fIpygNGxd9yCberKsZch/L
qf/MVhGkU3eBJUX/p5piMj1ku1EddMgQI4Eo974WniCDg5HLFfZSgU/szNTfOfCi
MHUqXMnCDZ5wqSFwUQFJbzsflDHR+kRYK1bCTQhPfiT4frj5tBSh6R/7SifmrGnh
5TPP/muGC7p2oSzTQmpuBbJlj8EMpFe5qUntFCTEeIn2luaIpO3ieCmy57/+QcfU
uQMZV4JADhVzH+s+Ob0hPr99TXKS6KBksWYIq84MUV36NvXoOjvCK7o+rXAHjGjU
ldjfd7UtmIjngQCOcCZdHaTwC1TOLOChb9xGBKyeAhAX6iMSwJFzW8TDueFRzizw
CdxJ4DYANfK8MZprzxzseBnR5rX4Y+IlYs9OGdljx82QdNb2ShPJSpZGAHCJppUP
oEaJVBjT7pbi8plCSrapnLFb1H8rznWcw9YOzVJ1EeAuxdTRF/avaM9IQRTWoXyi
zc9q7hNqokB7Vn24ubX/4DXBWDKa/qtFfweFSsHx+IzX2co6BifohcaYfFSGxBfm
6/BS3lxwS25lOzhIa9GtNVnVwsSPi7ssWbEKjizn2WLxXp+RcDGvfHG+Kw6SfQ+v
Jbb2L5kH5W6eYq+AbD+TsZb19xk+UP2vzNCjuOKhUkX+124bJdAz7PFAKDLzqFXn
X/sItjLKnlsCCa2oaUEJGcPAHji77hiQs1Q0ODyD5w5Eh2LtRgW4VdLzC2zuhnoQ
ciq1Hl4+36y+FaoLw05V6QqyhcMl9o+JuwOBWGXpttLGlUQxl34wAYaa5DgKYcKc
GJ9kAX3dragpE5/brM9EML8HPoC0rl2eGxHdW8jHpjjycFzNLyeA/ha6+4+M1mQ3
RC4iyJASPNAW3btD2fsMQcoSpqGfqCwGAFDK5C3Rg2yUsTn2nXaMF8NyZDjZKW0A
J8jf7Hiw4SOO8/uSIi9NS0ZYyZAOfoe5STsR8BuSgaoq90gVth+UiNw0JmxJaUGV
65IIJjRRV6s/9VkvbBsxPlMtYJsIA/GqCyuPtVZ0IoWLewXf49K9Uct7uWrmZD56
teRqfwLPmc0/upu2Idp224poTdNYIqf4w6izBZILpIK9tL/4lZkBGMyXPcqEsqAU
FGm+rkLcqWCn58fbQi8jt2rQxm93ZRwYUcGg+DWyikHFbOogBFya9MKLwtTuhK3J
BGqhEa/34UPoEVVkQdU1JuzJv7Pji+rPquBR9qO3w59l20Tw//6X9zwKN5xNx9Qq
7QlNs/XO7G3asKkZrUjBLm1Xv+i/OxDgpXe9Lf/Jz8z20SltDC5wQTnFNttTn8TK
FfkVT9SzNiYyS0WsjEdTj95ZLcLUE9Ju8136nLwKAhdlpokNEfeL+ozffWATyXSO
+2c0FHjh5WfOxQ7wEuMrQgeulqET2CWybnny5uOzMQv5eqgxujAI5e3t2C7LCbcJ
G9y1U7lizlCBOTDU9UJ7GnZmEQ38he78EEO+miw+ylOmQARgTAIN7BDuFa/E1gGE
uJzc5aX7rqQoSY2Ssr2A8DV07VhSsVM5NNAi+Se04znlgnD0N3RToMFNXnNI0oKb
IjOGSTL9+f+fGClrMiwVtehkot++m5GoMvgosDf2ZIctNlQAhfP0/fKUZC8QFeX9
arKk2DZS9kdkSbY80zBZqCJ63oVuMwh81mWRXThUbnIEvG/APSoBXyWducgZfrwR
Kw2KBQC3CHQciDyuYodWr+8WArLMOFonxMerDHbzAVVKb8HGqd4Vd1vXkH3m/Zkp
1KjUy/oE7d0ENaQBGQNuNKqDbnnsoyP076DDTwOVT6vCQ/YjLp7KjkpUKtQwZN9d
0NuB3NVxd4Qi+0BGkocvGGg0cPtsER2GLlCpmzT5HxtgjVyfftfgwkC0vuUqJ5TG
tsoYynM8GdDL/bVUCuqQI8luTd94fVFxpdYmxoroQPIVRnuYig/Dvw8ZuBqKwqQ3
wWCmNd1YmOuDAqvIJY5/ibwJXCJLhFwCejL9/dVkwapZfBBtJ369SBzdipm/72MV
EkHlnd55SucfV8Z02DB+RNcy5p39+Ng1+KrDZ7mGkrWFtXwMfTo4xbf3LlYtdwiQ
rWQnH1HWEWNfKQRh4u7hm4Htahp9H91M5fBK7RK4+KMhDOdecLfu7f468j3tChUj
Fe54LwRTc4wzbt4Qp5kmdyYFQcUd8unJRqHkqcU32B6QwNwgCD4qGiBg5nrwuBkF
3uqDboak0MbxO1b2MkBtRhCA2yfGhZy/L/KPRFLcI5Bqr7x9psYKoWbv1uajOWLD
U6YBU0FUlc0U2HQrXQpB8eMj9h99WQL+UIBotGPxZX9kPa4e1TaAgkil64JUIB39
rMlcBKH3wzqDMuqVLrEcOACj0LfuDT4DvQBjI6KxYhAGf2Qy5nCBw6xfuySvbg4l
u3M9Jry/C/ARdC9NrvWbUVkof7erW2VaFaa4uZzqvbk/zl/kKR95J1ix3bAVxK0C
BTRlCN2+apl8l10rxeVo/7WWBFBqaGZzi88QRamBcbIKLiWxr7JUn24oCZ8Xyo68
EjIVKrjZAQAC1VvRGPI1qx3ehuU95LJW1wOLPIOknN3/zSnBVssmTsD8XfFDhGLS
EdpfUFYveA+tnaEecWI27m3/EguqpekN5+jM8X63Puk2IXrS5ukkEjkbps7F6ieo
dQSlMrcFq0Rv73c13q/bHUKDBMBUzXgIfWO+W11oOGGFZzzZbeVIQUIJre02NQ/m
m23Ds3tOrbdoc9hl/sixy/ywgGUadE8DrE+cCBPJLp3SODFsLvblTIDkYxEj7SnE
KQrkIQwPsoB2Lh6b79WfFPlzypNYtyRVOszX8HyfyxIwyqOaEGXpt3hExLlQ0oHx
3cdxKLiRWL+hPBJkokoKlzMydpDtKxU5Z9PrgSLHFW+FMdZTDwUqEdgpgm5blz2f
jaKWYBXSq1KxvjHBTAFjHjebibewSyakGkcU2BHfu0O8pn+pqhQl1X6rFCqHNi+4
EZRWAyC7bVzhbxnNWL7U5hGRY1ulwmBpCEgTwhGnV44ter57Ef0HgxORjWcto4WQ
rldSmLDYycjkSiA3Na823YXok5wPYohfzaXT4co0DmC0C4yr8/437LC6lGenuOom
tlssu6RH8FGLbAmf9TIz93lJ5Mg5uYRDrurJ7aB9CaU4nC9rGWJr/uwb/ABHgw81
pKzZgWcY5FO5LOGG+G81VoTEntKDo/7MV8YMlamVN7X6gUdR99NmscGF+uomLXJC
CXNce6vyn/Dp9//d8xBYiUf0+zjz19Z/DtO+SdNhDEMgFcCNmNigh1coec+joMOX
dZYwvAaqWelgRk8egPZbz5gC1aGPVsLIw3vvQvOnKkCKHVx4lvfDxf/M3ATcfcip
Iu6EJI5lMBxItbD6yamqeVituO43/zEnwagrIqkvOEkPvzjPeiQYkMQCMrGGzjk0
ErEfNkfqrDumBvmK18hG+Ry6RmbPw+iCZfF9GU0vCcZP8ifyuSIlOlhnBhF/a5NQ
9S0VhreIi74SaiEKMACHNoS9Xn0bW5nIWctr5vhhKaosWep3Vh1A3O76R1K5srda
L8N68+8HsmiIOL8RmK1ju/9FxKi68aJuhUN9bxdMd6sSitubf9yEiGLARm6oG/Pm
pHXcX/URuRK/Pc0i+RH0YGSk2FWnFiIteXyCdcaAQo8EvUp7MKvAjywalZA92ziq
ibClGLGnKA2qZR8A3/SKLyJGJDphq2t8pCjNxY36+jZlniCsQN208nEAGwkurJcS
/grvKyEBz/mWvGpISDkJdm8T4qEfh80LR2KBsYGOpCzFPHubh44I7PSrY9Yrl9vd
wICD+dF2fg5baIjTKrPZXppWYysjRYXHfJxvi4DHlA+3jl+qqGLwuyypCQpfxv5y
qswOZyHtw1w3uZk2eCvZgYPX4Im5RaHt9X7WxTH3XovCRNEE/sa0NUWghd2QSztR
C4GvQJgXr0XHoR6Dkie5ooS0ipQIYs2qjBPWB1xmdZiExx/A+hzzn2HPnSn5GOWl
E3XnuJvoo2DMxCoTPa9fraHX0crJNNRb4FoxKfH7l+p1TEYZAj5wyMa3HP36X8/g
t0EjAlyXAeUsy0gVcFeBCu/+wlRNTQDjAEs4N2RYvk5eEweEi8xqnyuWAnBTeRUs
yy5niGXjYQCYW9zTUyWaGqYtqEgWWBEltmj0oplIn04dBF4zaDmVHfytbjyfMSnJ
CUzw28N/68ehEldRD8Rp6GbmdHW/eAy0xzryTic5OmPRUYKBhIOtJt2Wou4OWffD
HmlHxloirClvpoMOFO5uGG4Fz+TFv8kOFu0F69+JJMA1ONstybX3Xk8+1y65O7Ey
i8OHXio4ChzHEKLs2BcE34kmhYfNMtRtN/PHczwxkXU0NcSl9stnsQ2T5TDB0R+g
ZvDJ+RWZFCQ4wcTjqrpTAQAP8/P+hC5QaBna/aw4+Z4YtNLL0Cv0I75LmyfD+d+R
JjlViHgMCbAtfzhSH2e5RC/VHPwqFJWwOlMjARScjH+DcW72FgGQEw81c+d1xaFY
BsPW3EpjJWez+tLA6RCnqGVnEunGW8YY6CS4uU+kg1/1CcS+2j0Y98waFX5QQ2b0
/yFgX9kiEARCsZZ/gbot2++HPab1tcddcq5Vpj9asZ4mtoYzkKlJi+K6BRBLqGuF
pS5LFStNDJqS7SyOPDqAxCR99DC7E+ezUcQTH6QmMW4peJU+lkHLf6ZsEh0nuRjX
T+6Pf18X3iAbazyjFJ+WF04jgBjWyuF6+ey82LBvpqq8eWg07UOv3oSQzWFAlpXE
x7+1XTmIclrN7GJu0LKorpvU28LYX+JQYPgJfn+tJy1TRLMqhKC4LuVKSsoBUe6U
njTB077ShEUs4rkmmciMmNpqu8QDFHHlKkU5SJG8cjRdP5CQo8UaAhhJJvecuqJW
lMCdLhH3BYrVyBefPTYwI3CPiaA0au08Hn+i287uLo+p7VkZtCRNe17cfs1u33JO
EUyw3qe83rgludSFFzlr6ohmp+O4MKW9+/99rDcrsM/PtSJCMMfcsINMlnl4K90J
2RoKuNdPF4bi99QxrsPNqFRJjhindnG3ySYJYOpz6mhJsDRKfpXTa+fs5yAneiQT
7+kIJz5DtzYJmT4KdZRlk3McM5PsWL+cmYVtuwyuS/dLg0lcWAh5nBmcKK7yZ5JW
r2mmhkZ4rzFg6HfzyUpVOg+04lmuj9vnivISHayDGFiOsVi2ngwPiMusWm0GqEFd
td6LB4hi0DBvOeP/r0UpL27UKn99vGOWStrCsfVb2wWNSGqBu06eVRa6aFVgwJUh
USW7j1cgfPW7Z9pFCrXF73MzBAyn2Okm8jkZDsQ4QXLzH53eSzqdu78rFVOvhLxo
BjN3t4B0fOreqUJUW7hhOLKo3QJy/59yW3fye271Q020z1H5C2dpkj7IUtVxkUiN
ki4cylcJct5ZAY7kut6M0SxfjrvgUaZESeRCr6M/SRYMD7zkBY3MTnuEA8f1j79H
zE8BaCClJFZpb/BDPlm+KPeuuJT8c2poif5tBwDk6LJOZhQ4aNbB6wAPzqUSbjk3
82To4AJKdO2zc72gyakkfnvwn3etO/WsG/qq18bxKABfiDzJwdGf9uSfmqYrTMkk
a8i+3w1anAm276vVF2GeYpXSwqBWj/qTUfvEAMKZto58As46oBlYXy8erEiZb/Fe
/zCDooomMmv9DDPyKgm9MbuvV8nBo6Lsc+NvVVS/Df1Pp73SY5c2FqRhTiyb1YpD
W97qlQIrT373N+nj0j8JyGjn7TpqcUo51oizthiOu8tQhvwAry9xMOPTKWanRHvs
Q4Jr83y+9CX4IMJwsj6DH9vvrdn1Uw2kgl3x0jNo7TXTQ28otTRr7ajhtT2ohjO2
Z7AXdGqMPZCWj/qfEFYC9IjKOrRhnRR0Oxy2VpEFzxO+wgguQ7J5lPHJFRGyJ5i+
Lh0JkIruzfvNu5mqRqcnaxgEjUsI7LV+6JwIA3cWJjHv2HwHtpbKCWpF4cfEH0+2
Kx+UwetMjeU5T3Oay0iX74yXlF1hM+W8meUgXprSUHxRxVrkWcBjNit3R/6mLcl4
171mrK6PhcM2TIs87lInysL4AB8SlArLF6ioMBq5mIFs8HP/kdTVYB0s0/XIG6fQ
EhzSFCoRXSS98DWx7kO8EBrjd+7G9m5ShyznhS5Qu9TNYYejuv7GFazyjVOzdQFn
2kXJJXViXAPMkTCXWqvsleR4IY0e6WUnEZxMyppwDq4MUjgxpT86NQC5vezHz+cm
T20xgmvJ43TKBtSh3I03xkqesurIa2dmgoyAxKXonM12IV2nHaJRjD13J6wmRLLH
YjcBsB7fSE9HPTKE11qw6J3R7Ey7oJiC+3AedAkVG0CiSxl6CQMYVXj8Fp1qh0Nr
vYgWzuQknstkFQJrRCTRcHLQb0c8hrdqc0uErP73f/oaCPRpqyBUosXYBUzkJ8a1
c4V5bWVAEkVj59m6posHSlf0/c7bfKk10sz1I710O1qQgapVB//PB/YBTPvViuGG
O1a2FXFnwPTlyP4PeOUMXozJDzv/LMiscaxEhpYeUxnDcNn3CzL7SGjRDshd9fDL
su5iuPp+9rLkD2HymOKcFcBwgf6UE9QzwDyqP9juK+52JDsJFQkzd9ZrXD0fokr+
FcQq99rooYmhfNsw8lBr1LOr2QGnvOK5SWcu59NwQT6kA0/1W8Q2raO6Asmr+iyf
wGOhl98kW69EoL9foeCMSYUZ2fLdKQCfHm3RQPtKHGZGjc0gMvWdKg0v7n2ZzcxK
wmnaZUgaUlrpjaipGABGJQ6O6hYuWXYQkoiEp6FXda7SxoR0IFlQKPOGw+LWQVlz
BFpupy6h5UiBh9SjyxwZDJBzBAj2ZySlK3h/v6n4n/UrcgCXPUM/1k5CzIQeP3yz
hl3/IisatbjbsVYnMjnCXNwBcm8awoHFsxWFbWDpGN+QYFK1iKTcV3rQxv5CI0tS
hxrauthB3Lx68AlhOG43c5IDkxSeFwPdlGT+YxVVoPjghJCLB9s5AKYjmvy6dFWi
AvG1u34HpyUlpn9hxPiGHevS3wsb9Xh0hLZL5hf3EYAjFSBY5mYxTW9mGrmeYvQy
NGukCnQPwuReHZKZIEADndbwYDDKZGG/3nGcv4EVyCRmbY8Z+XX2KX+l4qqsac4m
/JFwHdWvXNLfy7XmpqZxXYDlQQmQ0V1y1MeiXrS0L7bnH1J8XyTl4aaXFFWyB0Ct
K8taVKByFVVgYKk2vASuue89vuzOmwqWIjlyr9UCYj9pbiXPg6gUW0/PjdbHiaQa
DqEfAtFfe54FpIeiPmwIAwscQWi2OacPsDAtmOFzvIIbaRmz1hML81W0ORAIjelV
wPYCe4BoFEi6VgGxmH0AY4ZxSyvq1ydEog8/1W1L1ESHeKLbpXiLIQgzm2JGDQY8
4EQF+3+PfGoivs4MBdeRaYXFdvaWGDIfJNKaI8iA0XEJqLq8ImiCUkaCVQnQ85Nm
ijZqDk5GJIM2eIo07zpUXHmY8fuBROjD78yay1G+RCOCF1ZLRmK4BrFPrqJAt1RT
9J/1wXB00g+r2qvYA3RKDt1QdIVliP1W4mCGJKIZiqDR4ad2cAroLtrIgre8ubr0
bs+eWcXngMZcDP3kRSxAaswiT/I25WSKyLl0wT2h8nYhBAFikIKNIN9vqGySFWwm
MZd/pmv3iaD1i7abzkje8bCJCDvkk+OAWuPwe6s7HwF3yUM1oLGwK832IYluFJsu
Dq1QdnJgwIwPtjpt4yBYrEGhWpNaAlAtL9ppm+KYnOZWoUSF+UzZtENstxz4Hv8K
ArfTYQmhwGkRonTP+q6YAuXXk8oJZUoHPM71LkUwEGfDQbvlzoSt+bPq3Z9Uf9Cg
+BmOsDoEv61HV/rTtvdO/SNl7HtigiDPwuia/Y5m9oMSHxSLvZrn6/hbeTys9Il3
kJxSNtFwhg6wOEsAey4kwZ/VDLp1k6pyU5iWu1640VkOSXXzY+8/5k5Wj5+AxYnk
m3Lu8pBWysgyPjGxjqc3qydUiMEmC6oaLinE0AY750YAhxnMgWwQ8ozKt89JR2WM
HdYuvX7PXDyZne1nbNrwgeZUrJBa/tWtjVVlxpv/EpIddPr6jveaa8Erz7JNawzQ
ValZUcj5bFgMoa3OatA6r7rjwngET1XeBXtXM7sJ+dUDy8gVdT4w4uw6xLpJtanQ
MzmpN7nCBDZPtDjO+sOKNgw+qrAqgVs8++RNsJYPPvmdcKOjuT3l4zRI20eFMmUc
Ik4COBcnlrmhLj7KFPHLcQSzwIn7Lc72TN5cULXczMorxmab5FvaqIRbBSufug7R
dTpP72hDjxZDO42clx8RKEKyfMrm79VKPI9fmmatBv1RFGlLBkOyRClfqJz5afiG
97tvhWltT10ERLCUpE6SrwsWQZm6CqGsYk+RlmCKN88SkB1H8/z8HJxtWxUvqUfn
cr7KHxPWcQ/tzXleIEoZYAqc1uzSl2CE0D4MgTfAP91AbIPQSUZvPDveG9u1PERX
RRKyHnJPhWP6DZnAAKELXD1jdtxe3GccTeuNRHuSAGFP9tvQUtmvtHZ2X0WWcp+L
hk/GWbQyWP72IAu3NHUGSUpgSYKThBUft46kVMqRw0A9Rw61zoKaVYVQAvhbsxrz
TRiVChex1Bt1HmaBjQnEsGhjHGGxwGcQ8HKStLri/vMydJtAmnrTMRKVUkvM9ZaI
kQRKy2KavCS/Kh04J3iSJaZVU8BElkgOdQF0SjKcsjUbRAPXA4r5b+q4OGDT+24A
/BvCQ5+gb0zbMgT6y152pPa7QD0BerZO8TwG1GBEOrSESGdV8vD7p5RDIDBileK1
B7zTwdiKY4EIw3NycZ5uSFZjMsCVDtK8YCAUREG4byC4LtR0/RDSjaUA0LuRy5DH
6/mGYcJTKjuru4Oby7mNrPkwvX6gnxeq4CmvUSX7aTLpUldTz0oBXWG+FdqFk0qn
JV4iDYHvVbVPzL51Vv933/L6tRCkWt8xjvzyosdokm7ZH+G7qEnLxgnMSpP3nbJN
3N1segYrSjLYGU3SVqA/iRWpFWCVqWIuJGpQHhZaTxg=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LJ8Pupvqis3gKemLEU+ZhU7z44qa3eYhmhTuPvklMXDR9a5lDD3a86g6Yz51Mek8
fQp8PW9H2zWf5FNsAr5UuiTI0v7uDpZIOnIu4VOnWRHiJ232wYgfNjoZkT58s/1z
trZTtG64It6r9SCiS+aoBc1ul3hXa7N6ZSbUXnQDbu8nNby4Y7iDf2mJauPb/yiK
IRLs/mxzc1HEHgb1U3FZKVOWPHbsuo5KcG/GCg6fUAAx86GaylKANs5Gje+42CiX
GLQilDgFkv6GOS2txnAA8PDevvf/5aNcdI9uYn8U5v1s8rTAeNFHYHmHPC/hpFSB
Pst+Yrbldxb1tP3rO0/NHA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10352 )
`pragma protect data_block
CfXazT2oZlGN9zcxHyweaNRxsfpTnuEnaehM58GWSPtbBN4unfRzCO4DTj/11cVs
mZL5Jph6bS5zZ4udbCAgNMylJRDnIazCaes0GtU0W8I7ieMuOWmblPDPbQpMpP/U
pbdZyuUIkjRJxUdc94LWbn3qQFVjeHhRiqhSY/Ot4eKg/OLhPmWWfhFYRh8va7cS
ggn98US9AL5qOcSka+Odgbse5BRVuS2cpytduXX82rSJCuJUf+Ny7jaGvjWQJE65
umgnKJIIaoLVQMxgBv2Pf7LqaqVx+0ihD7RRpIPtRt1sPrYgodHUM6kEUMu6D893
isR+6FkXWgKZXEjW8f7WmriI2ry/tSDhb+U2wVK2pRb4Pv1ClxrZHQYJ6F7tqIfq
nbXW9tlFVOrLAQRg03Y/KCCnoJ7LS1vx23KsJNDb81mdYwKH9hEsAXtu+E60kmxg
QZIt6gelGhwq50guoeccAyxP83T6tiAg6/9OYBItz4MsUa4od2DrcPfG4JIq74Vn
65AemzB/k7xTN2ZKZejsCuXlfdmAn18Qq3IEJxIS31pPg04Pjv6OHNwrn+lQnwQH
uIlFHMWN3pEMrdOCnENTsxDNlnWD66dMQYJjtCQapL8X4M5b5Br978dtg82BbJe3
Flvx2N9O0sLcveh+3l6ncWjVTabENfq44QbPBOfn5xMAURpRALb1JY4Jv8Kk2S2z
RjsjL/XjtdJRQD8qCDP1aa9CXIiE/ha9c/D6tHSTKqKQVsyP3jaZfKQlDDI94UVr
RWgK8dH2iEIQ3BfjQ3mXQtN/oCaZhWchRBeQAhsjguII+XXMIarX4MEsNrakSlun
JATbZ9bnehzwJtXKQYpYkOPW5SGgCnEdH8jZx9r8wCrkV8qwRGxRnKqrxJ9cs5H2
t3xUceN1xocibp0gFNUWH1EPY5DL70TjXSLCAkePHFT+GP82D3z2Wc9JVjoyUjb3
qPTnOR2xTocQ1JY+/K2sGzzQ2y2iVf41OB1oN96qgqTL2vPQrXy0Ndd7XnElAEVw
63cyLb5OY2rHlXefQ87aweCvzQr87SPU8zLEPw2E9aU8Pj0k57tmI64kCQwxnnCT
tEHg6YSKmpNdwaMnZfv7elYPkEUtnV2IvX89wwpXlD/lr6L0JEcUBVGk4B5X6i+8
oOUGD2KJK5xNJRmBRPK3wkXuVD0HGwBWCuxmbVWhyvnrPyZnRumxJFG8xwb3rxbx
ePExZ0I0VyhVdWh4fjqiRF16qkBPX1Y3/9XDADS2XOMA1jNVwoMYq2Q/iR6Tn5tO
fUjZq1I+sls9k7Yy48jm/fxp2lzH/NJmr0e8BOO0xbcKXxvNEf+HhZp7zhljPnFa
aRZskQphHyQUxYnIiZli57xIZgjHGr2LJHuBDXLqRyBFwpNOxcG/eAu5eFs8nHwQ
LqnWIEbFDX4uQMV7mrNmUfyb4UXUlpTLw0j9N0r8H3fQZlqYSviWBiFr8Qbwcrhd
3foB/14r527M7rA4KLpCU3RoVD4vkEkixIv6zHIRtj6kQhYRTndkqRLQH7wUHb0R
dCj1ooX7rs5UcoVkzSC4B6dN99OLQxOKUB5RYTA2Vnu45fc8GTMFeok+i0Kr5oVc
gmssi/IzACkentruOj3bShI35DLeUMU6q3i+zYuhH4GGRfiPp6m2Yd3v0800soPQ
KOSiOSbE9FzbDTmANId2N/tUBahFS1v2vRcqJ2FfMpzGYXlOu3gTiS8Fv25ipPte
wbNB+BUP+h7XGUD6V4ELwipfsKAOgb7JjpiyvrExe1hLuFsvSlIZg8qd/Ok+y/D/
b/RlhB42dErFqorVZ85YA01EE4AFqF3pHwNHVty5cwbuhhTjOeW3rhVhIWern3KJ
m5sz8+HOzdLexc5ritbc++z5bFKdVLp1xT2XSz7FBHnth8Kk0MSGiqyZ60CpLltq
g3aiMlubt9FX12fysgLwI3PzCLYyAY3DJat7cC0mV12TIciMDSoqMprd2SwpnXcG
3livK3w0OfioFJCAOrR7J19zNKyfDexKztZA6k96LjrMQH1vwEKlz6tVU9/2mbJz
jBIfCo0K8KfrPgBL3L0nKh+U1bhRZLjYM9Ydiz5NEPs5VMrvLXTX8ur/cVXLtIgN
6ZYEv2Tq4v4nJ6NUAI1+QDkoQDaucpZaWmpfPQcbJsW0mGcACK9lcUEpQNRSawYE
cbsLhTYmTW4y0hHssu+hstF4aVG93jvwBl2QbF7LlBlovoAI1jXVKTkA1KLEMHL4
UzbEVdpbu9I7sWD5B2IH9gf42LZ3dsUGx0/AjUmRzGAPyxqh82t2vfspU4luzKwE
x5e0uamqOJBbPqJAvEP9S80Nt4AyWI+H1JVXvyzn3BxTt9MumFyELz6pT7Y1y3NV
mQYD3sjXhdmB/Qn9qwwEbSZDYc5htoFkDQKDnRUUKqBTII8vdY1iEbmHVZYSbfy/
sIaTjvfYdZF2sd392nzhLYFMoipsng5XtSHpK3cwYoE1vtne9p2v8IyJl0XXOPjp
7wSWQDD+DtwIXw+ZEOibXclxcKbXGCpIP6C6v4/JfM0z4lFVvWR6BRQi0f/O1iK2
0MMdphz108zWVdbCkzs46ZSPNEGpuB5U4s0WYTMJ9RBVTrrtHuj5/rJQePSB+oVF
7fv7IuMzOZEEfX74atGylAvG75MQ8X8YDiXpk5KLEK4aOagPuX+TnGhjCXrFqzrA
Yarfr6ZqUZmxg0ceptXTOnjGiq0XHTKZTfI3MozFQ2nZF+EvqUdBbsnq8e27IsjD
hiQ/fEFFFJFRzng9jiFF6UnoPqofmLC6o+ogCP46IBQYZsbH+a8zLk4RhLGkqo/v
E8phjRE1dxgZmvFItvhywPR2xRVo+/kuG2iJo0m0eH+SquFcUknMXS8VLaRd/0of
zXieVp0C/ZmKigJs5mnIFBDSZsydhOwKck3L6ncHaLyr3xAh/wKjvi6GHuIj2SkS
iIQQW9K7ma44JEVGEPT+aUQPqOw/moKTnjZzJdWvUfr/PIBeOImizRU0xPzlL4lR
xe4yG/ravsbUqRkZn8UXSYphBaZU5tiIj65QhPP/UAiwx5HK92p/1iBmMFGwkxBh
Uw9zFTd+MP3szm/zWZhhz+A6iMQPPs950y+gfcN7ZxkaUrT+5A5/rkmT1Una1i89
FO0vFPtHMq3otYRj7OWer0MP0MKp112F0yFTgAI1GE7s09Hp1nfmNKylrLFcQ64Q
pkh820psi5vQfUP14eQbxMH5VIubEm0sfxssnopzz79R9/jsJNZU4gImMa69o8dw
t0Zl5m8RkQPVs2O1uRUGR9Ja3wyYaWas3Y0OhbjZni2F2zohqrbg3q4SdWuHu4xx
Aa1dNtpby3tQLb+mlCu5H3wZ+FYHRTEpWm221xxKc5VdLGH0WOULSU0WOtGPDisr
QuF0K4V9BFvlqu7EU39fo0DuzPTy31USol1Hz2EUxeAvxzcPAcohKi84yqRFxTuR
Z4O3nLl9fBby2jQCd5uII8jVDnaNL+1SosFdM3lvdHYgdG6+E89j41rA5r2Tw+L5
lHZ7c4cMW8fHmwN2fnH1OYDxRn1RV0QybsV/c3pdIrutD+3a4i7i3i3WC/AD7Niu
666Pn3aTOPLOSqmvqCGQNuUp4EzG/mR8YshHk7y+FIb/RCcJS8ljg2u4U4wUHeyP
j/pA5+rq2eeeboCWz/RPV7AOuWUZ21rhk1ZQQ8zA4AXC6+9RnoOAJALJSnanXlXB
n2AZ9XUBY/d6y3iYe+vvxNPcsiVA7dE7vemlM8CU79blDatxDyMjx144rfOHD49i
u5sO4O1Lp5e5uyeewYchdfi6LYR2Keu3GVpzXkDQoQzK3KRTrWgcV8H2Kiso6gy2
yqPob+nND7p7V0mvrTmBBTOdMF0vyaQeu/xpc8LPTQC1SVq5nZoefhTk5VshKHHy
jm0H4pk/Dmq4POOawDhqY/oWPuB/Rxph4Qz8KXRb7cjB/vgIQ3RxghmFIxjICBjn
L7YxqVaE5/z/wXYQKiZJPrkIfUBTo8lBaXzbJzhTkWVmeRAfA+fNkwZcXD0Rxci2
JDcb4XJ5DdpvQqRvHo2KI0TFZb4sYvGE+Ofr+jtGOXFFkdY8ha9FhQMyqlzY35Lv
DqgkB9AuXo13b8Xwwh/coJ1exdY1R6EPse0WsFL3GzqAtQKHD7nmQHIN6R1mbRp9
PvnKrR7NtBI/kxIQTUJ01UMG2mv25TewYk385ydkAszGqheeB7BnKUDz4SwWxHiI
gmyBe5jqgVk0pFUK8r8SkWvV4gymt+43xNccVYiVZ1Mh2rrN5/1aa9y73pRkB+FZ
5QNzw9qYFpP03r0mRZp9S6N0axOcai3eMr4XzItlL+Rk3uD4NVe813dkJ98wFZ9z
WwxmpVJS7ZU7ittdXYTLthGCfcO7TOoqdBXr9FpwJ8YSuUvKRXbwOgNNkLmg1vWp
xLFpXOiYXLjAEQhXVi4P18MsugDgFl8hywv4XsokkZaVQVk9vESNumRGeJ/s4Vaw
WwbhCXjHwnTXkq/5gxvh9g5AUHs32thBlMXGO4XnCgOzmNPWyfJvZQAMyYybN33s
xUBKH8+H8R4ewiuh+tSKHFZkq7Hqii3TgMZMx5QGw/9pxWBnTZC+pO4SY0LHcZC3
rW3kd4Sh88QHr2j8iiX4SBtzS3GOdi9K5GFW5JPsovR6uhgzoBLK+ZqzTrtRACtA
mMtZDXjRvUQ9HbTyGvTJBOmd4B9TnY6aoZHnkRzMtojdLgTlLqc/+33bl4zXF1+c
cgMRGlagPJ2kxOHAVeQU51tKQdaL8FIQpxhB2BzBTIAuhDTN7fLTh8GN9prTHG33
zhCyfLeHmlpM4JJuBoUeJbwmMXhA5m841hPCrwt07b//lOUKB1hvQKkR4rcPPvYU
uE4NtaNlg/TDOSXCEf3yibnAGVI+S8QsEgu/XBM21XyzilD4hF2wHWO/etH6tGy9
ZC3N0L3WtZrRxSMJdmboZrMZXxjvXKh59nF9w9fvhh8n8/zKOQE/Jx83Sf15x4C+
9QmLiSahWvGJNwQJYssAHBqoUUrta6Kp+Ef75PNLRszsspR03FumOYNW7FhWl0G+
xqXuxBIFuTK71JJ4X+YHJ9KO0gaEutU5J7xfUNDGfOf/LhZEW2Tik5RaqQRvz4di
LOhXSLkoAB+sXt4OG/t2r2LYl+xxj5yCx5B63u4NmtCVdbppoqoeWaFjjEguT6rt
gymYJ7p4HU1TmMD0GW0gZIzmXjTwOI065D0FGXLui/LYFosHjweC90E9WM03Fkce
w3nSHuLSHh88lyrSD0DYg5sTIUc4NltVVonJPsrWP2MYJakTzzf8gHWwpHfD2tjG
KLUjUTNJTFJeR9vJi25b+WBHCAjRfqDrtXZuQW+PxygLF2i7AQCyIeI8D/T/Z6gC
22dDr611rC7DFn1zMYWiq8Syby4ajQDYhqjNxtMLswtgHA586AreHdJWPsRXcC7D
fSBLO8u4QxYtql7o0qFoeF002/o2TyoE3vuBcDLKaIIKHbhlCx2VC4F/w9V3l2Po
dE6O9W7VjRTIf9t2q5crE1RjhMqgBI77DbigqfaRekwDoibU92FGIO3wO/O6+oZX
sEgeYNMNMNQ5q0kV1ucyYZubICbyJnv+vl97pvm475J+GxeKsGrc38MACJOWo13u
Fk1OoIjYK7vz79azFR6kKRnzULHNoREd1yJpsid0MD06xPBJyK4/cj45frldaOqQ
CO7OU7G2LdY6a7YFvCJysg1xr9edvftd5oWANwGJLSAcmqTMKT3xwFN2hZfwDDAZ
y+48zN1RR24nUN428uJQBAik+VUiTQknUM1mdu/3rgusCQR9jvXkzMLAeiuDUmTM
GIc14rjPX+756UJZWjd0DMzl8tuP3Nukeybw3CeVYsAhPvvXRqFw80hj9dcZmJkJ
h3jK3yojHcD11EiSsLo15caiCoDPTe1A7ZlNvqr2NojA4sQIbNIEX8LD/TqMPFFC
MBt6dEzQzHa0qlnxBMEn3s6G78a5aMbnmeme+Gb6aqIh1dYfSDNRW10BPEiWq+Y0
lI4QyrBVxWmzaPCjM7EmJKcHKewuReT3yomVCxloNh1hlgHT0jykwHzeiKdd//HN
WHkp6akBMX6fd/0UlxrCaj7UUWX6EUHhMKUSTl68ACEBq4BpMRsRJUsdNXYKQytE
q98BzQ5HUq4L4hhkOSX3ORvXk7kqaLMireRz25g+xUJWnSi951oI6Z+VfcR7/KcN
8bjLXlLNUPIl2TDMTRvf5FPhcCkO8t9Pj0xfUoAnT23wDKpsfFLEMu5ZvWvLMujk
uDY7s+KKqLF+aRJcUxtfK2KQATo7Xd1rTHYeEAJY1C9Mmk0S7DqkTIIAfuxI+JU9
iYUB6uUQ4stHBH8Di0caW9ubEMzk7bYRvM9dUuDn5lb7LxydMISQyEU/RRx8EWEM
eF0X+fg3lrOkrhoJugEHV+N5NKeaXZ5akStm4bt3KewaaT5GKz8dkIKsjEIIwCWz
D7Qy9hqCossKOzyGwRwkG9fpb5U01s/CDs9UIHoXwWR/HXiKYi2VVcVi8f7Oma4j
zepN2sTKyYE+M6MJq6zwigsPufq5UwLibeH0PGNv7BIflUMYvkVzey/yJTks2iZ+
tE5etKh8XhYqs0p/ayNCTIo9ns5Ew5MjgzXx6INPBz3SFAeCZUHxsh4tpTCEKHum
BJs8j5g6RqFgLjz5a3iz9aNOvVEtY8FODcYK2SDDl94mg5tzothFLNsfX7Q5BQJf
rXQpTsgWnFbB6pzVvsDv4HA5imRs8rAVeBrAJODewCYTTlltB4s899seBsfCayV9
W0j93NZFDRvqy8uGhmlS0bRLW4CTioJBlE2rnt303ChpUes4rWUDIRMOA0dUgdfh
a549JnO5P82ex8uC00qan1ZDXfGCz3LS2XplJ+2mrYID0NSYdhnRLgL2OGs7wrj0
Mhe1mhyM5U7IIhiPKPIeg18rVi1e/47Bst5AHv2JmXJEncUniJa5lbvRKArB15oB
3dUBPUa3QxLuCyh7O4I7hy6NTyW/u1oIeTu2kbmIYsHU/h7cxIJzHsgYxeDGbgJv
5igjrIyrbTt9czIry2Su8qwOwusdC52ol3/h6x5UJ5N2/CiYwt9AeQUFEkOZf/0U
uZWTrs3rZU6ORiec2IM00vn2jbOPUNpGRJnFxU/HYUZAv00mWmRs7ImSkfZydZGj
88qcaNxkVH9piL7j0Cx2M7Stnzh5WUwAb9sqr9WJ5Cuk9RLc+6GGSFLNhcwhih9L
GZYkeMFalZA/dJTLwc2kEpDkE35UUI0KtroIRh1oVp6cNFnx2Sgm7Bt+Za1khfwm
qCblVrhH9IvE8nM7uARhHWUYVcqJKgibN04qjpubgQjN2qOxxnH3kQdT6WiBi0Xj
OdGtzJnfJJ60xXHjXnmOUuc8mQXmavz6fJGvPFFh3g48ImNIzgmfetQ6V5bXWNz6
4mjc8J3cLoPJSL4EzFfqyVfxQSSMwOIj/xq4JHWd8HXkTBmHI9LJt8QhMUcvpRsh
i79ZYxb74y0MwL0GqTHJx02BYusJkByW7hF6Z3uNhs2Bur6aS7AxIhvtIiht3+27
80KTFEqKAnjJwVgagnaSAiAdOZFFUM40DhlIu8x+v/JjmxlhBtIE7O31iH0mwZWM
SYkO+9E7QkHlIpo92xnMZa12eesGG2BN5cxiX0iXsbT+odM32Nmqn5/emky5oGTE
T+jEtt7+qOHwU05gtUElOpk/ZkVJokHNgXgxvaMGkCzMNGc32E3w9O4hjcFQT479
Kv8VT2SjvVX3Ig8tV6zwhp/mBLQ9zavj2053GvGgr6SK0CHiXe8sVFXtm1iYextu
2/FDzbLW1Qw5Ls3xyV1RMlypWu+3PQf1XdK2kziXxAaCj5QaIPNp31EppEEEEUvZ
ubYjhDstRlH3zBz7c6NSujdZ+0fECq0EuMjaMZkIu0m2lHzKffKZpHPc8wUa7c/3
kgileKAxaCBHdNDrfJ8+2XnqikhKYUervj5tV1VDLwy52QVH/yTxSbg/4U5KrvhC
SbWHKzzKnlKfP6kWALl3cf//zjkQpecV7CqyQMVKSNSSn9iiPv87jmIZJC0O1c2K
zEd4Jzx1pfKLEz4Cak5N5rFIAiUkLwLd6A5qMRMAbIfpPQ2TNMZYr2bn3LZToWOB
MjSgerkpdBXzq9BGaObKxIHBtq0hukwaEAVw7E4f0dbdmeqtTVTqDpceqoFM+xes
N/qaSrZMFuPSFJGlyLbm2KeyyWNqfhSYz2IcwvjgWxFfL45up2LbksaRSIN4uQHa
aK+sT77rc8NsRHnXEQXk+/8PxDp7DVhaIKuBP2Nvynjta7Vg1vNLTPoT7S7FUaEw
AnSaznio8gSkAYYsdd/2n/EBp/OyYIoZg1iJx7f2jiG1cIneRrK0YmCgXvGdRrIe
OMQjMBSYh7tLZjBQxux3B9k8aW7O45XEv3WtdwL1Q2DsmbfZlZH9KX1Ndph9/U3u
BDTEnpJSNl0+aiDbjevLgF0U18hPWRNC9e2BHE5LzkHe/bgoGG0cYuCLAoytDKYe
pXXPvd+nD2a8RtniyJSw9EGTMuRUu8B1rfjdXaQwLraDM3w6R3tPvoOyZeserHXp
miJrJDfU3/n+PCs4brfnMM+Gr/ubfKTj+PJ6vdo7mp/k/fqBlPOSacp14Ivaz4I1
MjfSn8dxXFsBYcA1zHN0YP+wBxtIS3wee3hTdztoXuKddSivDYIfQ88Mfk8m4hBL
e24r5kgmuFUBxDGzay3Io3CwmvEtXvmOb/2InxcFYRkJE8ST7yQGZUI8UjXS8+d/
X+Y5xpO6wpww6vLqHue869iPm30M2lx4n+5JZJgB/33VfN7OYz1Nkjj0eRKGU8Tn
SeU4PhdwAjwo5NBvPVJZxUaAvl+vLHCyG97VhuqtJsEDFkW7FMxCkKJOGIJ3WbuK
pW4PX/NNsc74LpwpmcG/6VfhMFG2ZQPVGBfK4Dwv04EFOC/4vpc+I8bRIZhR45oW
U6BAYKxr+vIfStNMnHAzgvCdT/z0MM/b2ImzEar0voQwtfi99HK21I0+erkn3fOO
N3lCanc2fH+Nr42O3gBdDWDI1H2w8Hh7dMsJx32uQIBsxLH+HTppmvDd9dugPCN3
UDnVbe36ByK9wx4w9XTJcomD1wQKUp+X9VBO2EXpUA/5erOBSc51k0zav8O0a81b
+j4EsYr0sCPgC3JyonWprNLTsU4pA7yFQVFo3r8T4PbzsHJ6+3tgVxzhxZ4JtcFt
E+GwrWjb9Q86Pa1eMlP4njau5MI71QMTgGGnCDefckhUmFeNiEwZvNPE9jWkU0j7
FDnSM1wlXKPAfsc0CVD/uWXuT+zr2KHuTtiqCVfovopkszwGBxgeopFrxjoYEYc8
kvErgy3vX8GIXwvLL1YAgFqnIgvFp+iO9ZxhomhBR2+t2Rs56qEu8P3xVjAJDRgy
r2p35Vs3nDnrqD/OVmV+JYlzu6PaACtY40VFA3/bXaeb+5NVRI0oCGS6ohhVCis8
AOwOq4UxQMKI20wwD76y2B6kk87wBaB+0dlgfB0WiuC7GCjPyLcrp3Oqm5i0Q81b
f4K5etPoZI4rIQIrRNXOIsoxnO4AoHvaKVUU0zKseqG660lEbXr95dy+RtlFsH9s
jtYPelf2qUs8YWI2VVKnzWJLvGxo1vmoF+tgO6LJquZMyyMt0rOShIxndePej07A
YhHCxQyhGfRZWJDfkl6aw2pf4MX62Y+Q0Z7dCU8APtdTkq7qGPRJJ9zszBa4pwj+
qrAbCAOmAd8/GmXY8p9hrk4zVZzoZZsGeq9Mo8osJksTIzyY/Q3Ymu6Ea/EoGaN6
qmUzhN14IQNOeVVsT68k6aZh63z/kHZusO1FndXXUNqnQDC9h9Ei89gbyN2a0cKt
rDdA7BnQA11Gzy88SUFqLPETz07A7kBNZZXJLkmAdhSKBKHjFhTYkk/q5gu61XRg
yyBuKgNeesS02bKsfPyGuv2L5Vjjuw7lcaaYkAsmpDI4KN/Z+baqL6NW12EKD1Cl
c0G7PmOiniKDbx+G5V+57OWWRi08CZSNsWXPZlacd55es3gHjIG/XBCK62fFpx+B
rhXewaIcpcjMmd7p3pbUiS2r34of31x6TBLTCao1Oh/ukju8GyDlbe1PfRCtlinZ
Optg2Rbx+8XQJ+LSh1J9JsPzNeedHTT5wOrTrJEpfFw2+hs9r/WOJ+I18Akv6LVM
y2nxUklMuysRguaB3V2bDziO48fbyFNLrPvGHoiDCqtTRE5xqAWWFq6KtUwCtsJw
WNjxXiutGocYwoqaVfzInCSWxulqfZnBK1kgd4pOw0FvMm9Yt8FdHmoSgSetHHr4
Ywqx3LSI6dpuNeMUp2w6wIBIkccugyAif6gvGnWDxzwPJYx5gNWGQFMHHQPWuTGJ
FAaqhh3RKycqUv3eSSX37Q3Jhhzs0zBSeI2WOBMlVxTR3ChFPLXTnDW8d8KanVYZ
oA3XIlXw3N6ofiXK+Lwhqn01pEP2yCbT656jRrDWcRhDEKUWEIgDDMd8jFuYsNjt
fwyyOOHpG4VKT7aJ4/QzwsEWJavTgPYGz6ssKTWTzDdwfi3hvkYSZtjxJUzHOvEU
ovjLAGQveoH/RYIUpeXa1yvWeB/6Nu2CVIMYqwsQjmzu3cJFpoSRzeJVBjVUUf8L
sVPi0X8AWsFuNOT6EGG84DU6j40m5etF/Anh1Q8GUoNEivN3LzOIuxMiC0a0wPfM
E2YL6F1LN3LmrlBdV5V525lWDdVWMQGwT+Hr+xNWGQ5DhfQJv0E7BkLIkFFvsygt
Rd4M0PYGmaqsiNBJmKloBel0vilUuaFfGl4fZi3TpE5PtxSuP5NWV3lpGwU0XLsC
HBazr24g1DN8OnDUPeipf7ohHQ9DOxTYhogSMoSRwcOUG/6LNc61wd42T4CEd5tY
u2BycHIDmO6k9RgO19b+XR107EQw5Ld1oOMY/+8K0T8jEYzi8ENWaZ2a/G5x5FOf
GOAS0xbolUi20bbCOjXSr78IFEzuetfhKnRqrh+Uo7Oyq9G7Q+VeP60Zpp+cz/ZX
/4ousOdOjluDbIXdeXpgZ+mY+uJ+aOyQ9EnDvqS9XZj76oTOXXgP4xyAeeAO2zNk
XDF7qiaxl7YUizPy+6ivhymge9QhYhmgPC7+jHEz7yus+s8dZRHxAOUXwx/PZIw+
gChRSAkZk9CYhcEc9zDY8/nd7uNu77tPLZFJ1yM8Ok3v8uaoIKo2ZIuEe66QDBOW
WNvoW0g/eqMgUls9EPo0zreetuXdaFwCa3VFv18RcXFwZpQl8HY50DdHiEzx5LNh
+9aUfbjLq7JKRUkKcPN50ZXWcVeMB/az2kxa3nTcGUWAjy+In+eszma9UDZHwmd/
G6pmHZVtsdgeEItQpS3KYFA1mftQc8YveoEsjV8zQQySZeuPNpcQ5XT/JIZp44Yr
UROdLyJ2Yt1Z9kdYvZbt5DTLg2rYvgqb0H/fMJpZddlhlAv6JSgub93LX/0Zxl53
KLmFKjAZpReMkp3yLf/oQFLYrEBYUI9hh19JKGyrVh/byh6rMmYqltlKQ2PfGdAq
uIpa4leU2+Jkqd/ZbbLZ7td1UWumJTeBKy/OeCMG1iPfeTbjppJ8mBogcS2A6Lth
rIEChxnqEnTXixlvQjEZl8TurnxI4v5nmb4KYCdA2T4xk0xwmchvxySeAf9902kA
nDSxBoHUb1dohMZmSpUJW+QhDVYIeF0OhaUh/BfGtFjGS+8TaSf2J/f23TVvzIQw
PJ+067vV7KbcwvVP4m7QNwMZzi/BoyeufGXoA0GFG1/u0dMAOtgplMpssOQHk6gF
kCx3jrkQFJwhD8SL+nv+2JP+ud0aTA5mI08yTWsZ6EEdIxBwOpQfTMuO+v3aALKD
mPt/KuaWtuPegYc3tPlaTIqa496qeXvg7mHhV3JsL+mgNW2/TXN32Ya5GQvDqLWu
LcyC6T4QbS4O/M5tZh7wxrhNfgxnYDiC96uvZeR6YhM+jjtgxKLwWM4CLBQao7wu
6Eos1hPVL5rBQjwmCZirv/FcnlJFYcMNQ97IyMv+CZudcBYsSkKKtXbrMR8kEHTM
qbn29Zjy6AR8gWSFsK9yDgXKIm4ylwz+G9V9DLu7owK7hSpurllbfSLMPSwBDfQ2
0JDuYIeHSR7sR3+MOiVX98DASo/scGkZ5qzLfHP+zUWOF4ES+DmTL48/OkxnqOpj
uDlFyB3DdYhpz9u9Pw93f6Hhqg9L23dHxJFt4BO7ZNWrMh1PVhIy2GEAHncWWJwm
DsJ8iJfqALW5FNpYNZzjedGBXhfrudMIZl7zhqQtRC+Isr1Y0yPhV708dY70Q4+w
hxRrGYFoqeSrf87FwVsNIh7t4fQJuIU5QV3+lkZUQD8Iz6yildgd4YsiHbLEQzFD
gAVGxWOdGQ6ScWxAtINaWDdppP3hsIW5bzSh/2oc7DiHh0ggoSAYYE2G+OpOze4V
dGG4j1H/1PNG6XdTm137AoxNW9xFYnPMSgXsnsX1iGhd3IZN4CTp32xxWKH42h/e
rrsleRirhB/KjmqGEYZ+ZzfvM3/vbegsm0G3j0Etkf5G3Ft3LZkULQC/pGw0BIKt
0Iw566ph9uEPKgYCz0KsjR+dI/Hfbx9hFNnxOyS8s1R9gqnNfOm8/6TP7m349u1s
YbjAg5TFUDC/0EqTZ46sPHD2CVYpd0WPvklftfYbrRdrHj6xTjA2e1l1CDvvgVGj
W+xg1pExPNlBMrQyzLwZE8Z19G//NyLHfl8sN03hfWv6YCoXg3Z9bIuOYVGUnIH5
7SK17maFLNDoBUTR8yFcfVAPXFGqp2pUI+yp4fq0bVitrv2XqzxqPTSIZCCN8YgH
H0nNlHE2l7e6tOZKKwxP3CKlTXfAu7tkOEIBx/UUBUpGDBo4PElVpH2F0PGEawPw
k7evZ/EutvVvRiDzzRvneBEAW+WmkEZQx5HA5+2BU1Qz9fBlUQcvEVxswLLopfcE
fy0ZcPwRF9/3803slVblsw5xWJUMPEsgjOWISwYjKb3yNT6z+2lAU17jaeKwlGgD
MlhMYdvVetzv3ieyw6/XFQbVwdr6/6QSVSBg17cAt4cCWeQis2LjKKEp21tVlncr
7GkN9K11CzT8UFeOacqShfQBWWYk2aO3wpbfVuxW8ZtXtFfRCBMi7v9TQGh0D972
+/6qMy/69epeH4Z9ceTJ/RniRuQgPm4NHVZtvaeGcNsAkg2QSorTRRwuEtmdCM1Z
QZgXwnglhQRbXQ6aVM9GqkCyjeelnrcWB1MbvKHE+snIeKrl88vNOoN3WNccltX0
eVNz3A8xNggefmQpFw6hYfKhHzKPHYSsCZzXrKaeViTsu0nBTR3Bgu/R32qMBsOl
WPAtW0wacSCtDZDkKGaWMbbUcvxM7AxCW30jSKofqpHJNrSDbPH5O8QkXJvXuoa1
RXKuoyc7LSSBZjw6mONNw71NFhUdegB35WRmiD7BG6MfYuEeAl/h35vBBHCbJvxV
DncxNccka/9mGifk2NaCGMAApcwW4no+qjI5I4oGVRipYcWF+LZQZrlHpVkzcaz1
hZFsOUDX37NbYq0xpURj+HVCXujZnm/JMTTZboB78pcvs1mfauh103i2kdngJlt9
Ezmg2mtfWJVyPkDMqVNMdB/MYnRsQJIZQBZDa8GHdAX9qTIKy4hR1abR49Gtd9HL
vWakpEGh51pvGo41NXhQmeyZHC/Ck/5dX00wbAC8ecvbQ1XMwDlo+blm1Z5J/1Hn
RavnaVcD+vrkhgjsampBHFzlz+uyrwGoSsVPcL3T/zbvSFzcEAT0DWArjy+xVg8x
6XbbtQE0dRe02ZUEDLdtnb9/o09ks5N5FOiVeFoQHgw=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
DvyJ083vAVYebTvmaYgUzNWs2Uq3XpeE5mZ8Arek+yZp1N0XydAhSnyINL6uI3tF
xEqAV8xYxGSlsDosAuUsPCnEKq+u3mwNLZtmeFW2+C9R6MOVBnQvuqQZuTymmeXZ
Br5TwxMU1ycUkQucCMjK0eByYiNI61rD6FXcqhTLxalC5BxIWd9/4Ud689wPbE1s
C6sKuAV6nhVWw4pRzbqPG/bW6cvIOjioGXiHOKQWeA3vAFhDT6dw4MSwZkDtd9wW
V86kGCrVlTI+rF4Sqw0Uuc5Jbs7zJMDDhIGi+7aiqFgjh01WWStsVBpdQ7P8suuY
a2XBtwUDS188qCbnB8d9qA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2512 )
`pragma protect data_block
XRxtDOCa6f1WdYVgT360s/JiSb2qOk36iYHkoNMJEewgd/7rp8BiPKJBAPzrukSM
UXZsH3mEEvfLQMta+NM6x7Z10/9d56Y9UZJzUU7lyeo1vvK4OlrPkaUeJK+1ZZoI
ov7DJmXWFVM6deV6wHrVf2zuUbr/Y8CH55UlowSjWKkbskpBR635FH0G5pPF397b
e2o/yUbEwyQ7fF/sWyzbf6FVFGadIqZcw6fgr0XGErMY3FFV3YiNvA/EmDRCHoBi
qibo17Fb2ODprrUHpFFSfgDTIBJHjZfI7UhIUh60dRgnVMRzguU6Mpq5qh81VMzN
Pz612hsecDImNzNZkj6+OVr6DWU78ZuEaAq6HfdQJs16Sc5Tz9sYenkdF4PIrR38
xMbARvaz3FGeyHNHEJbm1k+aVyogAuYk85KczEl3DR4HwFsKDvGvhPUEV9/h5tJd
p1+9mKmLetOCqeBCj7djub0k6qmV5g62lXVGADw8AgPqrgefbY2Mb+yKIt9hVMMk
UvyP1Ouiuvy1lEt+Gm0R0WXwpF07ww0qZQgGoqbmcbDAxyqToL/u8SDAbOsfbOxE
iY9zEcPKywVnj/OtbZew4fzHeg12jNVFx6VWvwvPvK7mIQkCCqWELeufZSXphjwS
a79+uFY2X37ZH2daD8ujN9Na6LMJd/bYLCvwJ9Sw6Dif14XbC+vGkIhaQ2YEiEju
swEMjwXVBm2/reCL8pogt4iPOjt2x8J8yIP/WcTKyQwcdM4BlKn7TG3dUVzcd+U9
Dw223OKlueduWcZi6FQfo1lc1Nc5dafLDLCbxZmiB2VLZqXuIL7gsb/ZDfukTpso
tR9bYEMsfo1EAQFxSj1AwebyPfvvYdQjvBlCMbdfxMfHHIdeXWvj5Fi0jhmDjVU8
3pxavmjsX34Wr/tlaX5ysrpUJCCyM8It18xqQ1NNuh1YWN32bB6As5LTv8KI7c0j
u+H9SV6qNB/Q+YVu5jQLG23ty3ykjkaU8w7x4Ru0m3eKESuJjuQ+/JRx64YQzmi4
ICsyYi8lF2AlrbUjuJGcrcZLjvRME4lF3ArdbkedAEhytwMJxSvwJj+SzlVr9yXf
HepB2tC/Qz03zv+gZQNeIycmqnBI5PWoE4vtKDsQU6gHJp17PjY09KV3uBR+pNX2
24TVFYoSqsHp//Gcgw9jSwcAv/fzbXFsGi6jU1TKfbx1mT/2zN0O328XiZIiR19K
ORw3QE5l6TklgdioTjauVyDDA2DpizF+UHDFpzxlo/6iraYV4HhjZqKf6yg8Qpl3
E0fSf+gxSYu96EqDsmPFDCJoMJidL7Gv2qpxK5GYbdlEiYneIC20ze9Tm+/WUohJ
L3zGXYSlTPfr4HADOa61sG+64gqWcFLyRSL7KpZ8GNtXzdOlkJdoetgkZ+LHnJMV
AWuQWN243ukBMtXTvgjatSJyiOwA1CcHZsMI6/SXVfD7yoJpw1TUeC3hGPa7T26w
7SqStWlVsy5LJlvMjj+3L2CMhKUeeFzns6pJjLot0mvXI755Cb/nQi0liEOlAEmM
E6YxEMvGAE6JtqpXVdxwe1cGC/8dT9KNLQXY3s41bjAO8wqMFQoKutVeYebCHWwa
JrDBX4ErnRHh28jQ7DbrtScjMuM9RvrMz6EH3JQ95QTxEYPoaFjnLmuS1IYBLSp+
7syIKvNuWwv0+qd2znz0c5BVLMWg/Z46H6P+EgKmIRhTF/zD8OBMJ00bWGHBZV0d
VxkN5b3zg7GPtWMl/hQEHmY+zJe/5qbYN5m8Wx2o8eXlzLfeoVrBiQdvtJLsy/lh
XdIfURzJ46XRZpPzkkb9ybtrnvW/14rZx/tS4tMsp5RFuyJiYMDcFISgsJpROcll
IY4fBVV8UxmF41zdRZV4z65fC6rA2LoigqG+I+uSC+pwprmyhG517xWHZiCV5ZOl
hVUNmx8E9dWVbRaXLbicFjUwbZIHZWAIv11XwWeslxIP+9lpeF8YNC196ik5BIN1
8ZL1wwljjkrq4evBey9PNz+LA99VWkwqAr08/dnLp4Da2ck8Wk0CZxa3t1phODNA
sw2QGDE6W5Z97bIH3ufkKndQIh9fpevqV4Y2fomT0vGpXJ57OJkdPAVaFK5FU5tU
NFyJdcuIO5ZURjyZB9J2Sf4TnXQ3Iyob7HPh0bx1bQRZYtIi1qNhHLfPmuh6+0Q2
u7L8ypo3E5PBoUtaM4ecG/yP5hlbiTtBOjvsEeL7bqQ/v+9QAgCCrC8qKVWZmvmO
HSC+KNw5x4Bg+hi2NNhLPEmb6qTEAtJHfq2F1iiFD+aqp9AxDTV+3HUywqYxAZNq
jLueAN0A8r/O37+2tJjRPHwr72EITeL84Yi71m5LRjf8dehk42nkCQWaZubd8D+m
eiMyM2Ord+0offh5n+5H3Zt1E3YUnGT+EfuE55c8aGCZPhbwDc1icrZREYJO4Sgo
GTIP20peh/Z96NxP43tHzMZ1vTpXQjLF8gQbLcfEO3SwYFVec3ga9VfPKojYVFua
UNCBXwZrRY4K+rFE4vD33VaK2FltuE0Cy3dF0djgKIlPn/AVeJMbZyC1Yi74Ge1o
/5GJCZgqzSc52W1lDRnu9RAxcTac1+2Wgbe6DAAkQqrOg4VJQugCTpxvG4sWmBOS
eqsNPhnWI/T8Vpb5+zhKfsy6adlIcWL+BfsLZEM/1eJGx56SPU8xVKicP+I+o1jc
zaCWcaDL0G26tjlc4rtJmRCouCjReZFw5GTJbMtlIL4NuJ2wqxzWcsKTRG4Y2f/l
CnHfDU4DQxyLHEM63aew8fKoQwLAw6yWvchSx90LfVYEK1hqeGPRdLVna7oIgIyM
NnDy2Ki88mFotEyEg5lzDTLG44/in6LvqkwZ/FAaw9tv67ODTa1rkjQD++dBwNUt
JCBNjXNUiT2wdl31XNKjNgEndnq3PqXX0gNncG9ljmoXExCwWaRItmIxJbQBqt6h
YzbvGex7WihHADgTpzm2xhTtXM87NC+Ki33vBF025g6NsGy+yc9dn5loJ5mijXGy
t4qh6ZZoxjDeVTyYTWT5eoM/zUaaJL3fD/S9es/3R5lUoF+pUo6C6mlTyLM7E/dB
aCKg3dNIlJ3MZlwoL0wu+c+9VCrEzo3a4mciaDVQ6yLwR2j2rTOybV1m/SUbo2hc
+jzGUdjdZOwMDjsmppz1vPF5WDeteZtMywxTDmiHJFrAlMM+y8toyQ0tirdRohvf
gFm0riijonWrZtcVUH6KAnZLdlJH6ZhE91fjcIQTPApmhorJez5kjLWg/DHMORVV
/KIZAOqY0DebRTqdF1Y6Ph3l0+foBa8z0UgkO1poRCrkcofGNuAY7ZitJG2Xyuw/
lyL60SibBsS8TSzV+7R1Qg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NZ7fpQc4t9Pj+XDtlTZaBmDPFmHLA0b8ld/xwkeFQeKdU5VzZFhU5pW7pkh+DZy8
URm+zBIa/AtrqU57ghFT8bJe4Ao1hfQ8yyjO6gIIQSLlDwHR8QThQXSARiE9k4Xh
QdISJ/aT5tFSQiSp5ZDVI1VontlmGprg4TlyJ+FCpiwJHIgqhGD+q2viVG/W3dvg
sYqYg5lNVlZj3fW60Ee/DQlrS003wWdbaShJdDilGWbcB8WvJJBQ60TEWWfF7X3H
MMPVSBhhH1/149rU8REEVm8NZqO+WitEDQLG3DKWjevBOKzCkVwZYj9wUEQ1xtOA
heXM0S+9XiLZ4tmXelsB9g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22672 )
`pragma protect data_block
6c5P6YuRnYAy6yzBe3qpT09NNg1ED7uVgDQ6vo5ONcjRutoIFe+EM28d/cqr5mDq
9pCHZu7RKNKiHkEt4r1fdXUEA8axqvNDBsCJUImfML8VZcpDe/SMB5ex0/CDFuHR
TdVpAb16/IaVAPsQmCeJeM66LKejmGGnZQ1BRRvUo109Reu3jguWODF105gI8SxV
KHINCH/QCjUSnIzHd2gi2uO0HGbU1L/c03t+YOELF3W+AJ4r9Wbzif0bVS1KKi7J
R7v/99Yz1pH2S4YFa7vMt3OTabN9oBfwlYdFTD8CleMbgfJRRqjphXFIh8EgCysn
JaCO8HXUgKVUCtYIeLyUzwALc37EA5YLSf7+eONY2GPDdnhMii7dYDVwaGTXXReC
R6WBITrhvbbX51z0ahYRgNh0QirmeLTRtEdrCC+Wou/DFJVNPEugafjkc5SP47tZ
AVMTbm7UrHTj9bPlCRhBWT+iTbEBi32maYqVLX4O8lk6XQvMv0cKmcRDgoT0TaQ7
cTQAkRS9yrIBIthE0lTPdlmQnCYc1fm//Kz93Odkrrrfh8q8xP3KRbSsNeCLCsty
dvQcPvKrf2WaiignbcVx+AvUK/BDmJn1OQvQYockbHCDyn1+2yhhTEnYaik9TqF1
tjaY6+sX2lpLVQHsv/9o1ehf/Iut2FA9iqfLxUBO0xurbJElDY/yMfPockbtG+rJ
V5OAkB758JA+0+OV/kercIScBGWJiMJYBJjCLDzodxzhHPi/EXXORsiMZvVC+LXH
U76+yr6eBMiB+TiNzxxHa9znwrsczzJzk1rsXsueDJnw8s3YGhcDc1WXi/kqbsDG
nz7TRzBAKR/AE54Nj2aujwnxJcjlqdxJud4VJMWMDz9BPAW3fK/Hpk96LqZ7jl7N
8/xgnH1jb7LK6oSt552AVdipIy8PzIoV/gB3UF9p6XU5Ku+f41hleJcaT5+YJ5Tr
GzbdUadpD3f8gTnTr4IAk/JXnDWkRkcOt6AHmAKjbA9vQnFmcx1r9kfGR9JhBxe9
+Aa83n2FFKzICdIZdOe8z7/DfpoP1ssgyKIl0t1X0lvwmCtYwvapSeKICnZAQfvB
3QLBUquh1ArLv0ZjeWCmdsHqEekZf/nUailtYaIcqSQr/WorGQJqDipYx0k1CZov
S5eIVxQNh+XM4v2FF57cRQ+PBzVhFj3ycvS0h2rLktmVQyzWqaCbU0V4njvwjA9r
VQSqFruX3T5qCHulLa+lj5aj9zlFdPxhQ8ZinMOKUY26vL8L6Myq0mlb/ArrzofK
7YAB+V1tVi/GiKVkFv9+peoiU0pk98z6E3pE/bM22NqAkgm/Jz9cT3plc1BTR472
sDLsolLS+oxl4gb6c4HRMgZea9xZjNzXmXn49EFuDg5Hx5aqmMKhCJw0dZ6hEWE+
nKBos1mGsgXZM1Mave5EwNpDU4I8aLMbUciWBchcuf7KKoCeCnCi1eJXu0QPQ/u6
8dXYHRZvWRTjwEEWGwWrOSLD4WxEvkdD42qMPxfcEjZUXaQPUqC+ETXmaQ1Uxm0Z
niWmBlPIQFbpTO9maK8ss0jRYhfLd3J6kElgzVyppMk0sH3+EVCy/Dowv4PUV5/t
T4CrhYEGg2ujLJVY+AMgW+PAHuBjYrYcsmH3cigM8voKVBuuBRA3jdTNAAtvLV38
K45SHhnNRXumi5DQpTRN6IWcgzXi5gLE09XDFC5a8LNg3rsLGfdlkPbqgEXkDvD/
2n9avtFpFmb0/ny4EzoSOdRnZFYpjpL9j5dfjSV/u8J3lPpWq1m5aR+vAIok3og0
AJcDYB0lZDpKbMQl30ar/m8ap1DG6fArSTd56nZL5W3oeqGaj4fswwtWkF7AYwtY
tPo72Ycbt7J8tySGpYQSuw4HIUVr3Q+VZJSmu4qFXVWLxLWI7ZYA/Pu1G2SDi9uk
pFZHNSUPt+r1r+/W/cr7c4fKV9vpQcA/oM/wv90o6/naiZohltcIJKlWQZuwlNwS
83wPd/SnFT4L+61SQ4R3BV0j6GIjpCsyMg5WKyJcyoRwIxw1mRnKEnI1mmU96+WU
LkoSfRBm4f3FruQRAZ/8iaTI+5QgBZw4nCjmghjJkFJWC7yzUDiG+7Y6+Kr/NJ5I
ehg0+v7kXYdTaZGB9LPuhZg8sTVHtauRXJAAfAo6bB3LBy/7QjAG73TDUSFLynjo
PL0RnQbCvVZMwJgqYLN+LgyNKGo/LGVbw0rDz+F7pHf7xpOqFpCvO7dGUPeni6pG
C+nIRZnJs/88IlNl35rAVCW+d+TFU5jidjNHtfGJxMx0cIUkn41KBr2N4X3y3sga
w6w8X96RzPE2OXLMRvXWoE4D5DzDhccR1EzpID1icUXi0IAax96NzQRM+LxzHMfU
OHG0YnWohdfn/ydTIk3AZ1TIHDrU+OcEl3vo4tXKJaY3SScSNhguvpSF2BD7soXu
As+jg/XOaaT+jpXPexNz9BmYsRFLKulRS8WQb6gegaQdUtN2tjCiLa9YUyLoIVJu
cabAgj9vn5BSBV7C5EU7pth01GuQbD+lcYDwmgiSWLeEygi6uNQhvUk/P/nwbGmt
KRSmY+4fOGLmeE6OWhrJnyeBoNzCsL9h9dPx6MxBg23w2zvKVfnlLh7yu7aFmsXQ
PY0ejw0fOUo96f4AM+vLGIFQd/j+dO3BwC6aW9rchujsAXLaMqkYF+owJ35if/AD
kEB9OTwAkXAYtQSTOghW11J6mJciN8UB6uRG2uJeRqI2J6w3YGEiOpYn6JMw7J1s
LW2q5ZMwdoWKuXHqVqJT0sZoQ9iiaOmW4jEmR/TKSBnAljjVUt+KAKr25Xr+BxQp
XDGJhCjWzUBdHSdx/6+JGnjQ5Ubvk/h/r5ECIP/Fj7E9GnIwqWMvjZktI1XTdRqE
rcs0sjvjSItszKVd/JJYZ/8XhGA8ei+qVX1ykf/Exr2B7AcTaFlg7ZspfqFj4Rfu
juYjmbNqttVR8Se+6wkO8oSan/Ee88FyWRKESduP1tAz5au7hKBakCeX3g3QkRci
tAEc2/uLHalIsLEfQtSZikLpl2+rlj8aO0emb14NEUZ+WFYdDJVzDmq6RYON2mTc
tYY/LVuAvhcRcpC31wunAGeiULXWtwSaq9zySf4z13EYFmdZLJ+i+wU2K1pldNBM
CIIAofTqXYL9FSFh8Anaps0PjEs0GCgiINNaqZBcLAV9tnxYIxlNDltVFbOnQdLP
ChtTR00oUJduBxMX6wexad7OGiW6klgCLAJEGrTJqLbRgwlBmDjooVPkIA7kSq0w
kwJS14cl4dupd8QxDo/pwxSpScoiz2kLo9OO0w5UdxMxCu4pzP67UtLF/ArdLfVo
2vnWifRZYfcW73NnXxz8112mKyzOMIbqEg+J9zD3hyKzcGXVmaJWv+Yjkng3iFus
HFUyAbjrw4buzKozAr7dY5GS6NhKiRKnsH5fiop8tOnstIXqhBawYyPjnj3cm2cK
eu7pHCxnbJ0CJy4IVQGdw856bR9UeMzz0j4QsE9UEIMYMQdGmIqqmQyoLgdy+sDz
GITin8mxf6K6RCcbIqtljk2o2CamiXehWFzkMjv5BjqQyZ9qLVuJpMz7a/Am6BUM
ypvKaPfNc9LRcII3mP3BndCP7pfv34ylWqN+AzlWAveicf6wkBYyIgSIqwreMbWE
KINLhkkCdt1toiuU/gWnYyCgQR4pvQrFg3ZhFKVnkklPrnxDmsJmF250TC03wcRK
4PETEqulgVOaOoU1TL1GCvs76hIuQnWT0hEf5awaaiOW9MSlwGO984b4rS8fCo9g
LwkSJGi1tXkN4uT+Ss5Jr7x3pmlz9dyJm+Ee7UWjX+5rHwNGji3ZKfgBua6eL4yP
FkZZKQLlYMi7nY6SCAV77VT3Km2LA3023rvD9tlEcLkMzhx3uPwgW8XubPQmUSp5
xZ73ItWgbO0Z9JDs6SqML62j8P8LwLOTEGz/ppJnkt/RNuKnCxggQEgzSDBbwnrD
QtvZhA7eP8JF9KJiLZbUuyHuBwVCiCmN/BDfA/FX5pbXKM0EkV58Gt/YhVoskEBw
4Y6dAA5IWCJFIVSvMG/pdpcSTG/FYEHxt0MSTO290EzyS0Mw6moD3gjoWRl65T1f
kLwqULPQV9ffoZngnNRA/Y9y9fk1fQJyeIInrtmmQIFTaXyDyBmdxv7Th+VmxEPB
tR8ei7L1pG11ZwWdFJ2Avr+gLaNdJX26QDg7DuC9Y5BxDaL+yw42eboy9ZsrXvnL
usz2NJ/tkbPXSAXI4XikwsvBfzib4+aHyrJ5/pX4cPzE4Jn1viEIymqVBabPe1aB
36EKE8CA9YIePcr2kbnnotpCvzOniW2a1hJPKCruV+7y8Fx7RFIOUssQfFtgLigN
m/xif1adf/DyEmrOEFU6gWNqUBB1ib6R0JqyeJnJlFxde8FNjIAhx3EoPfWk3lz4
xLAZ8OFYF/ur5IwPASdMknJQUOTJ7RbiIpihOTSkuDA2NT8KvOB9GetzspW4vhHr
4ayohlw4mp8ZFcqCcOOJVBuyk85hP1wDGkrp+eMdOQo0v3hn9djE7x9Zx7JDKjz3
5cuhmOIofz12fRFXDmROvURnsfAbQrg7jcOAWJWT//lDAixBhmr+mEvxk7H3k1dV
hKedpO4ekW9+dI3f4k0DB0TKN8fyeXfPVRoTiqNm4A1iNDgLveQH6ua72wsGSemH
FBb7s2B+VPSXrU48/xXoePzMh98GZU7l3znUXPHAChGCuMuEkTeSSEPLhZ3THae4
07IHZNL4QxgIArR/119LrocDWnnPOYKSjIis5gOfQgPS/OgSJAtb8uVxcZfT/Tqq
Cab+lg4LxRoYE9mkqoxBEXdqr4lIDS5sFIH9SMIMbqTiSjpQZs5JZLIEfeGgZH7/
nSivXlayJ44YTGm5C6eGVlx/u6vY/6zrMooUTCj6AtBtb8aZbQp1L3q2tFdGb+mP
8sdnjCNjKgCy8j1sH2fqAkkQWmYh7SC+SoLi+Gw8VAVF3xfyCQrCkgGH9Myz0rJq
VhhM2dlRusQxOLsFETuH12fX4mQlDnSA6mVYN+q2DPp0CTnt3e+BGUWM7EXwn+a1
gx9QZGmr2ztwXgfJXAYu36UXECJcVD1xaBgxqlGh00w0fVfXpmVAGVQLglvfWJaq
vG9CjjHkFbiELt2bXGSuLBhoTW2RWRqjdw8D/zuHi+ZToLlD81yYvswT9ec6fmoV
RHwMhEidZVuminQzoo3TblSvRIIQapVznwB9nzXtO/y0g4oscYkVRODHKwxp0i1Q
ObpFYViRyc7iLUtW6838WPc0KYCqSZ/N5wJnAJjpWWq0sIeK6pITy97Kbj/rNvD2
8IrMWQDJ56DEjkbPBeIcj8p9RKV0fmE3vRB+mbSyHuEzvktXBHMB9Gdp87XTn6xz
Gx7DJvHA5vunvFnCpFzWThtb5AN2yNJsKNXqhIUkqpdcuqmActow9uiBRrQN+3cz
SwKoFVDT4NFKeyGDyyfcC8dAbqH4x0nN4BXKvLvQnXGnTLDDXLjr2lhdq4vRk1Y0
dwk9K6B3KbrV5LeW4NTC3fvh0syAEH9G+jjt5BL2GY+BuCouKwL1PdaP1XUycbud
+WGok6IUEo2YF19Yz4sS7AOT1Ply2zKgB9ZrBi6Ksy1J1h3R27vZF0tiF9LsfpST
PJV0dtQEYCHEY9xKBavEdMP9d9nVf95JsZLwx/BRkJfTx5gV1tQd6vF4urKsAXdI
alGYdYyYURAToCGMRRgIRbv+A6QnptC5OM5os5MkdfREo70z+0ZUSf0QtExQq4zH
3zRO/Y4WdtMEHkPfHVtkrTLL3T9q6PPJMrm1OZKgQ5QmgUXmm1lYhV2ebAfRkUm4
4rUjR900sNO9qpYBfiShHaVjPjK9Wx33RPnW9RJ/koj7+iQOlolskpdX/4jgWHHz
k0THpDM8Plgph/ua1YTnzlk+3Dp83My6FotgBIUiURXSBMViaLZD1SE7pxv8LTKd
HT1VT75zLzl7/RUCj+1GYvgq56z9XHJNeHayDto7bXBJ0MzJc3CFLPHkI6PWsG+/
G0ho//lqPv0kVkIu314q6NiFAtDnfoffRKMl295yUxZVgYpkhoGTbKBNmYBs6iLx
VY0bFu/1Qof5t9rMJ6spWcfPJvgaW7YqA1PErFebRv9PCTj3zIb7ytht2Wgtwvtj
JllsDBO05iL6A5ocuWzWPbwNKN0DtTO6YyEsTeLB7pMN1JkH/VZFI/PUbcSgtTOo
f2UifS5kmbnjsWyqXKsORAP4QiZk0PQMPnlirl4XNz56JzCNQsQ0Lhmu4DMqHnoD
7BbWu0xOrPJlMu53mm7q4Pgr8+7v+9DRbrA+okBmqEFHJ6N2zwaReaBuq12K+7/F
4snu/PhhilopOCFd3CwY4gYjRsjImZrAjgJWjlu1Ql50wMM5CcAyK4Y9M3yXa0wd
RywTXrfN2SEm0KVEP5QCfYGCWaIXM5kQZKkrduRQ8QImzQ9jUlsLzfcvK2zmM1nP
X8PyY+9F/vNzPzHnxxvdOFpzhKCUYQIRZSLBbmKtpqRL/lxSzC7/q43/Z9ZF7EN3
x66lpHP+5HYUlYyX+52+yHMnJTe80Kgo37gsHhUDj2P1voetS5YeUFj+EqeEwMG9
ON/zYvyofcRQZDfodhbT7lY61lZi/IojWl4jNmzn5KCw/pbXbW4171jcdxbJImSa
9LjBDfjEHM2VkjMd9sHpidnysmIN4/momAStiiR0nDkY4d5O+aGcs/GHko1uYCsj
LyikHUW/2TV56uf40S3frreN1KjnunV1yjRX4GpNJPD1YqJYiNwjry0T3oSW2AQ3
bD4hAIsqhYuuMSfd4FFf69hVVSqlUGgi1AKm09+D6CF9/sEJF6Tyt2CfdVrGj1o/
n87fY0yLFjHbXGqW7UguFsnY9NoRLmZd5HvlnU1hou4Hh01dN4QNlO4kTh1wgZUu
2ZiM9LrE0VoEV73Pss8QtLTubDyWHEUUgmlBhu6VULnYe4Q3jqQLoLbXBCEfAprZ
xlLEUy3m1SXk7B36Y6IqC9CwJujuHDyvSuqL2fJhOelwKLlyHrMeMg9WvRXXkWiA
nVbpBrbsRG2tSVvTUlc67Dg81cD5KEjan/lGie/15qkVU4cN2nk2F+N/DNn+/1y2
whMIvlvDWYn75VUzFZ+X3RpaQ9Pl1zUieno3xAxbY3r18U7rx/spHhLkVCdLs89g
aKSCIsLeoAddq91T/2xYik1j8HF3dGeh2ILAU+MZz30h/XPfk2DM5iqQRu2lPg+/
8EVmuBGb0QMXiQ7F3ZrCSoaLT7otJHwgXSkKzqI9IR7I7unaXByZvaAlpV1179WH
uzaY2E5ulEHseTdnyunloIkaejyGelCPf4eaR+/Pv7EJiQZqjBvUQhgIZPTbmaaR
wpiXRRlXLpkUuDnM3QAevHpljpytozmxkraqRTfZWcYcsnH/BtJYtKGyIq3bgu0e
FGXQqlazD7mRhqkNSHBT4RsG61eEdOtQK7fz3mWrADjjKX2akYsipL6EWsljje8e
s+WkU5YUGY05aq9iFd+ELAWrhh08bAwaj0nZTTJpx1G5QzRamGBgrpKrlXCqf4xt
ORz5nQ2d0+WHyMYLewWo50TEVORL4BMlpYMr2scKOA/nbSTsiuhyJww0uMb0jIuK
nmzBrPKvAxYY547611hpfsiaYI+AKaYMSECu5ha+2cGvSi2jcomZHZQPDXpJRHo1
9T74Iw+3yNlcnSOF3lJCNyubrWLnopthPPJ4Pr27Qk4XoF8vZ/RRaCIzFStSOZMi
oEwjl0NNPzsdmgdz0T+Q6Nn5Ruuylot48Qb5AhVwJRM5eDJ5x6ZY24TkiPOIVNqw
jz5yRBKC9jERKi5lGlNHaNjuUhg+kldqjZjGAFue7Uo4LwYc7ZV4yqTqQ47KZNcC
lvGKSK2PMOdMn0/crMPXUsxj3I2yvTJQn5PqfbCChh9a6DBNVmRjT6jmcJXoh0Lh
8jkQFdcz3VJ94r/rbc8L8LYclVZpHtokTUkutg80VjWW6pPZkOKDmBOuUXKwasq/
1TZX4UJKcePORRhrRyNX/0XGFtfzxYB9K/Pvg3zvgtZ0TX/KquMYEnFt8ZuyuK60
TcHik7J5vamtv1ywm5QNKAurVbsZP2jvldEpT89qbJPgbII2oXmomb/6jr9r1RiZ
weigjVxxSAlRivXjIXAFAX0JbfnoITYJouKbv6YfOIycMYDSztMMafoZVlDGE4fK
fPdvnXWIRnMP/kM4jfJOwv09Q9gM2AuqFoCJ0NOAnrL9wg+E/iZPcDq5xNoOEaUC
KKaJ5+TdDzrCEBNXmrdd1srlaWgfoxLRg2Zs/7uWGqq6xjnwR8Of0qp/bDwq0etD
3NOEihr08SMi4du8WsWllPnMDeN473srQwvTGGwnbOkBNG1Lovhro0nZah07MMut
QOkNADHAin3PLwpmJa1tfgsobBBM1ISWN3e5Z0g4rLjXI/Mhpi4fYQOIKDvIxaav
P/wSscXjrJdhVhIAdHzpHUx1nDu3JJVOMoZWX9GjAx/DPNsrIBBEgtnbhIDZ9pDn
Zt9fy4ut4nukDWwi6qxJvF/17csETfV4i88O7wuB5EXJiXv6/GQeACwgFx7Lcl+0
klR83aZ+zxjO31s+w433kFFg6xUVVhkZM8jCIJegVysTR7BoUg5n8goMKz3VKl50
FBiGHTxUH6tyGHv7W+2ZfyOVu04zlhJNUtYCRMaAh1r7kvYAPrMsTJpdKSbKeMCh
re1M7677WXsJSbx3Vfmx1pmDhpkwGWVcvzNsFmqGK4NOlhbSWoMuWmWE/ufbMjYX
n5rqLNESRrhdzPVqL/gmHLmZTY8YgR7wpDaBmFzdBeCySIfv/1Gx1LPRVecV5D01
B5PD6gaRNhcLMnuNreFh9PRxy+Dl+r+FfwAU7R7gU7CGPkpJ77A4X5sNyeiUmEUK
pHvvSXQklPcnFrBNg3GU4PS15gYiGpAvZlUHYKRg1xx0ReTPzIDNuMsBKGYtl3s1
a7lGiT9GNl6gLZcEphtvSv/VfalVniYVCKd/kKB8HwetUBCaazlu7FLQUfva7wxl
wrZ0KvP4z0tt3dtdpZ5WdCi4P+BDEArBb1c9NHdaFCuASCrmgMlC9DJMlReLkRXp
ky55Pj+KX2bgv+mI7g7VKLVWC/L5cpNC6vNqsGOBG/4orkoeKtcle2Jd/wBQi399
GtiRaxisrdBv0Mivh5AjnAPAkGN4hqCEJ/qz8Qa/Ts0bD8/yR9VQvH0YsWHRv/yD
MoHIFek8c/z+h8r9bX8raNYvPBA2pUJ/ad5UsMTqM2oGOaQzUGA5qIR79A78121T
mPWpri7B1M8wTCY57Tp0YpW5hivLCa8Er7IKsSP/SfWVi80c412Ju45rRGdg3+Q3
q3BH1d8mr0fZE6mOpY8rnWTTRnGouNx2HvT9QvZ7T0vATM2rXrK0zmhRvYIx8tzr
ODWxkmjpPn++5JA6KWdiQWwHefcG4C5kSFEIDnFMTpeAM5VBSD3fTIn6mCNFQRJB
mJqyLcZZPU79paxnyeQNSh861BgnTKvhiHzeg554/fcHa+EXq9B53WVLnOFAcQxD
bJ1uU/M7e3tM3o5Rhkj8oNkeYBr13pz8J2XakR6LDhrN0E64oaD65TmkHrqpsdaK
IugUmkUEnzz07k/H37WULa65BPYXLi7PtqiSRef7+D/QjWF5gUIOLff9OJJGMhCa
E/TyHKzEbPDOLOKgP6YWen5QBFegx3pYz4FCx0AmgTH2vZFMdjSFHoXynH3fPiuy
iTgiLxjNV7kgDHplWjOgNl6ldigI+yj/lwZoAa/GI0iUJW+RHQtAlP2F3RMyrKLv
mWOXClYRXwMQ5TbCGtME2obpTyazY+klXseP47tCJE3jdAIGJtLSBW+WewevyZWS
CDt3LyDiaJEdDf3k1Qg5pcUH6GyzHxVzirJbXAI66JnFKtsaANPbtFxFl5mnATv0
uXMF0VY7TEIzLhbBrfLiIkM/HdzCX6dQQXYkl4gUNTfu17NtmxBPJTt2R6CHwTBb
ceAe70+ii7AI7su49tD9iGdoOBR8/9ae8JMq0MCmt4sNnUx2RBHPHGvz0e6UG8Xg
5QxIOcZFpFcc8R2akSZ/Gfi/t6HyIOqpofAhjJJ0+rVxpoFdkKchj2IM/LvXz8Ng
9Aw/ONe4svVP1enYR7huCIqHwUb4X2sp58WpEVb9OqyynbWbsrUSgNecgkKwkqhc
f+v+cYc5gwZWxAOPDtaOARmqk7atiNYKkgGTbg9fxg5jiH/a9xqN2Opa1vubZZg5
7uA7plCWwKcUB8xIiaFVxPetwdASrWiigFcwTrSJpU7kj71n456HCWiN3oZiOFZd
MAd63ItIzm7kALQ51IsKhlU+Q/XS6Lh9j31pSeVlJQWLYj21+7/gk8PvnjhX/CbH
UJhsNzNQ4ye9fqcWe1YOkxSuaH2U/cn1LZZOQR+iCtvtLkZHiQcTu2Ji1MuNIolJ
LZup4ryWino+gLGWRJ1wOvL7WvgQbT2YdhqR09TfLoHV8fjsQK2ud6OR4GILsGCG
bqvOxFEczefshDYWHdLUxsBsC7YOa4T3ItPBAA4oIE+xBQ8ysrf1yZEgixBVkjtl
MoWSAjBFE+AjFeQgdKrjBvtW8/zfOrlT+5f4AoBlFysyYt2C9qeASBYd7GeNQaaV
0am5Rfay5oG0RTcuXTCEvVfe8Joal8uN28Mj6/oKp2ajC8gBps8goWWca6be18GG
UFAQQ43O+Xih+QFmy2CQA36SNzfIve9+UM5qxl+wgJoX/+nLUugviDriHLiD/fCw
QdQOWe2mulDnJJMJb+5CZM96jMiu0jSvD+VaJk5vOJbpuVkulrvTrbfzSqBDg/hO
d+KGj9djwrDnxSdCGQ4N9j1ln7IGqR/BtUDka0jtWZUfHmD2CTXEgx3SyGlJssMj
qqQ9c4OPsVgSnWkjKnAiZgvvTBtu2c9JL4NFIWf/7oxpUQcnaU7WEd/q/sSDeN3N
VbJnxEDpejSwUMGgPlSjmyyt19QElZ9tdshN5Kb64MbIHMDqTSqcgKO6l1RfGYmT
AMqTY7L/5Os0xvGfoPq90LxG3Pv6DYuKo2P4a/tYK6wewUv9pWLzGi7ep+qRujdt
eO+jFMqne2hcMpocVkH5eERBIuduynA4VoNnNMVzsTJnf4u3yyp3vAUTVhnQ7kTy
JmMaPkXhch4Mur1OWnUW4PJf9MGbiEkv7dkFP97nPmQfuD1HBb2Z7Z8S3xd+qlg7
AXu6HybHwbliZ3nHyFMZ0KryzhH6o06b8IQTp7PUdWjIWtahMZLjzI0lbPuPqvEx
2aMPXMMjC6fH0mw7r2A1VfOV8V3aL1+TOSaFro+fsp5raEjTVGwxbPic9rnYfjOL
1jg4G2ho31VwzjM6NBnjgBDZQXr3KKOSodyrjoaxQuHXSLO/RzoFuDlbO0GZ33cK
eZ/qraSOxbYHAg1WUA6b6t15/skD71CRYXyy1bSDLBHYZe8msttA2EedM8CPGWPO
Jfnb1f59l8sxOBz/Zq3dh2AZOAeh7XN8OytihtP9zho6UvWAV1t1ijKoqhSVTak0
0LunNO/02l9i7IpGiVLy2ORbJ9h+XBKrXaDiDN59eVNMg+DQJirQI9L7cnNQszpT
WhrEN/kJB0H2c/zJNhCe/eKbRxLeqHjLMSqOFH++rxzzFR41GUBlmrw5CsiEYJlr
9LkDu3rldt6UjFjqwOsCKzgwXplumD/angaZgmsTtEPAg90sy/O8nf2yg6HOy2P4
kGP9l7ZkDRWBj3hezR0tUMR+k9aod37U8duyjI9JAksnFXTQwgfHJXh93RzStNbs
1+SVJVEMUw5bguWWfyqX2BRou+SUcJQKS8VxwdGyn2n4kaHaboVOt+0ARBfeD7PP
+ALFchmpM88RUKKJ693t+l7EGPYqm1jYGxyyMsh08X7ddZ2FRpfi6U1vD3m9GJGA
LSZDVVvNHgUTRdb4KdFqb862AKgg9ID7X57VZbo514RqYr747Gf6F3CqBuI6pt89
okMkCxkQXJhIitZL2rpyFalGJeI1XF++1xU34wdvERqD/bcEuaoIKnSrp1kruJ5W
qivgF3Gh/bYmcIoBSz5DfeSfobMd3YDjBSDCabwRbXhucvhXl3RbOZWTtGouXUzQ
wU0sDxEVxAWWGEXYucWH3Bqwd/xF+JlmM9wCoYIJuJBWhkW6bBViCcrw/VltmUZ/
r1VbUTQaNruQBeWjWZ1cJJaB18W/Okrihr+EqyEYTrq+ZxvRsKm8J8ZwMEFb2ZHt
C1dBvVfBzdFROsywr44cvc9+k//ucE6wqhLYTkUzoNeQsyTSv3osbCAILZacjMT8
BcmN+NjeqOjMmHjx6ogUctWpdlWZRqzsj553SACJ65eZyFy50uIETJCZUhbaP5LB
jA+zjNswnfOfIgVi2uHNbpi5gtRJthQqWm1GO4rHWHIDRICbuqtUzDG7Z7aKUl6E
D8UwqChVOAGCkUSgzpcOCl3QXt+dmDWHGBoVAFIhb6O4iSYbsMd5TaBhcljY2kOc
MfyJd2AZlg1/rP2KxJ/2lKWnfKe3V/c6O1MtcktQjIo4CIcXvv/CUfCGKXWz71rk
nVejZgKOHrZ0W2ewCn9GvZJzY9xP5lvyaRDM48O027dKaGEWuN6DPHg3LYHgNOQU
h4IZRvCVpIiELUf23qD/OWKiGXh3BlBEukmlPGrTfB5JTo/NeXl4DgAUkVYBmpLa
rRJ3Et1UQ6b/mUUyge3ape+G/yd2rVF8x0A7tGdd81h3KrWwCaB2ob4nWvCxmwIl
xvtrHIKsy25gpXb8ENPW4Fc6JDJ8c3LiptGIW6BlnxumFioYtnwUJ8h8kXPx/geh
sFO2hRXwJpJqns9yjpWoBA4UQhP3nxkTzkfz1Ffk7kcyCLD/ZaZoktC1X62Ei0a1
fftLuhJOtSm+PCvcx6Yrk+QiOSYBRUPwSU35B1hiCZBRqP4IyFd0/pl08mgfEFl/
5nVCutTpBOobmRYxduq7ldG0wZpUL9egbRyOXIZGQeDAilQo6/f4FLmCRG5EzP4C
UqpLd+7OvHbe3Ho4D2b5r8cJCf7zCWa4nfwBsKSCsU+KDhlNNgeU5Fl8C++caXog
XY6t4lnVHY3bJNHSLrLf6E7YE0MCj/SYUuqe7Cn9KVms0Gl1DeRSZhDWtJOL/W9+
nRn4mnJXmjL/gxvXcHVC+WladMyIh+0rkJIIAKvJZmRxSc0xOKIQg8xdUsNs6XdX
TZ+NJXBnykbQmgI2kZhZFumpR1Z3D+J6ndp5vd714aLhwXQpWpyeyeFv04YtyaEn
Cx9y4tzh5WOaECYvJWAoWAaebeHc+N903+GC0k9EOF86fUO3/CT2lzbujkBLfrzQ
Upfuh6lGmdYfK4DJnCZ3dgHwDrMqx9+jRH47Ozh7R8UfJv41ioRCavZImcMMdD7s
hshrqsq9Hv6vM79y1XZvX3WQ1L8OQLx0eiynf/P1TE9yc46aHtNNpTth8G78zB6H
LgVjk3ARJJzWXoG64u0asDl9G+1QpYF/K/rOSBFC5NpOhE3Z8pgEWpC6JHXUK90H
rp6Bg9E5EO6Fgim1FTH0OMwScKph51CLGV6sYyww1WNK4218Gqm5dCi9isI8GBl7
7kBmazFhJnBbkTmVJXwFR2FH3fHJGflVupA4oQ3NZOsz0VUmM13v5AvadFt/18PG
N+TvRGHWWMsA+N0ONjk0bRWm8GqPNvJ+Fi4+DJT3TmNmaiU1WuUsdgRV11QHOhsD
utcOIDhqmU3XTusq5Jm4DLoMUbKMOBo6sD4LRokE3+QS2PbA2CVospJczF2iMjKL
XtNjzNsK1sx4m9ayYHykkqyHkQowMpiWG5eOGhhy7i560Ld0zCBJ3uoYHRniY0vm
e2uNownRrigXB5y9YkAIHkLJ64v8EeIrXktDxLNKvw+ySXTiku8x/9MoakeX71Yh
nh/7OnYCi7L/ZmR63kyXSm/hY/IzFpBczVYR/g+IogbRVK9QOXBI9s1LaIfMOdGW
jS4adnuM4J7+sb5MqCANXYtpHx183Rsh0WgI0FY8Ujb0AQyRZVfgDvNguFzSoLsn
0NWqYABAiPofcyqYLUiCvmQss41aMj39SgW04KyM7rLbE4v0lA+/szx9wjg3F+r9
dXtD5KHHLB5nq1d/oAWpYb8ajIbvwd7nQt+/PIsmz3JSVg9IIdvB0im4C+ijzYrk
PCCmTP62agkfdiMchqZbMmjt6Y5xYXSOP2XNVydEomoy+gBnlaKwv6gqrBPfq6mi
6UMFXWCcdy8fYQb/nM1zlMdhvbIV7F0tNtibwjyIpj+HDLMmavIlU6jo/2BOFU2A
NpoRD4PyrLSNaz7l7AEH25ma4rXwiUDZq4rbePp/kKAhNFuU/pdMcOQQ2k8f7vGd
WHZgFU26btej7XzknSQQdM/Ry2EZDT325d3pp7lQYjdd9h43jfO3sY90L2NFZYCM
/WMaQcE8og1aZJhSigHasU4xPYFk0s/JU20YU9tfzRs46fXDJPfjeTf6VICr06Wg
6+Mcuu3AQy/LFr6w2pv0d2raEgX/pEHDHQej2zucZYiuQ7QVroX7KRFx+lotBQjd
m5oEHDWDBFjZX6K8QhWMFu+S87ByaYQd4CFN0G6V6/BkUoHjQUjoGNEqRbd1zyiN
2wQS6RqnTgW6vgJXaYvAttzA51C1OkDLBTZ9CxV9EV62xEFqemRlmQ9fJ2Py+9dw
rYdQXtbtSLdqKdxdal7VsMvqZHDamJcpgR5DKq7qk+bRIMdmpy4vUvj5KsyG9Iis
EmNfaJNwm4Xl86mU820MQ0bWIbLGUFYWP9rVbEm8fCFpJzcaSpdL3EETcojJinC+
EScPwzlR8IggUWEyPEjESfECfIDCO1AX2trq+dy7D7zOUryGIV+Zqy1T+31p0uik
nUAsTBBXb1uuOLqXiyDG26iQS/xE9Y1ed70I2omansgrUYX69WPY6JtV8LNCKHQE
RDGKYoBSfO3OQfbajCYdQc3MXAJf0Q26KqDilZ9+6FrhAZtHqFCq43ZthZApPShJ
vp6ljidzhggO3sEAmPDUvfC49XO7U1IrSVvr7cbZGIx2xQsRtexn7cZAoEpa7vIX
0f36rXk88JYcI48zk0g/ceJG6YJEMOKzZv/DVsk9pBwFw3a3J9cvIWF8DWMKpg2v
eB7P2z7nymxO/x7Kg0+nZTGQ5LlMHrcrDHzTEWjacZlIaNqnLJoDtc8DYHvXj06h
Qu2vsPtJ/fKnn9tE3vtNj8puujA0FPWZn3v17cn/uSHm+ILLdn1JV4oyCVkexxI3
HBMd1c21yKHpEg/PkQeXUphcnGsYFsmqMTFbfJtNWcWPIALQXUDSvnjo8Lab2MHo
w/zSsMRrW5rdCTQ6mt2+LBL+HeaBCLoSM6PjE0Dk04FjL2Mfjn8C4GndqCrfzm5i
FBApNxRY5OuLgjHq/EZLvQ+L7aM18eKee/CAtYSdrDGXSixZ8AJldBWZeJJvrPdi
hYXRSTeI7za35p6NmL3iVVwV/Fa8HYfUmLvyG8NZ7LawE14R88QLcuAAMzzUXcLL
Nrm8jwoA7XMJ7DxvwGYF2rX9Nl1tjax6f2IJByYYeDy/G+bAED9TwEM8LJIiDLT1
b58ADgH3oPlLTqCaxJNDOhZgYI832mDLMx/I7zcTcdAC68TgmDk/aXZCtmdue/gd
YB2YT47hzOgGIorZbJPx+VNYZRWnnb5mP/K/NcE/zVP9BtYFYBvmyntT87sv16fn
ZS7kd4/go39Ay/SwqHHBrxCs2nzJqBTWgCmpWsaOuC96844U2Ovu97csJgVufjhM
GwU1Q71rvEliebUp+fzR7TCKHgKkeoJom0QEHJuy5m2i7DUFXLys9qg4LNxr+HuY
1nex9NriNk7dw0SI3UNcAUKcLtMcyJYTSQEnjYvBsoT2wOmxT+1HYKPZaJXwQgC5
3Z50kHdbyVQ7EMZbPP706bjAc+KxFjcdQpevZSN5rlIeuwE4VPy2s/QTyIIIK1RF
Wx6Hk1IA32ICSchRLXax0ypFF5PSkeGqa9Yf1pvTqCHXNWcBPDINmtiP5MDdE8FW
TrZn4X+oT/q52lvIbceu5ULG+yPbsDDuq96LSkJo1bMma4SjWH7ZPfA74x+pFfLm
IfOyGuc8gNWa/zKNQFW1c/B0mTJJfePiMXCak1aayZVYwechmqOFEwGfM2OUbwnG
ewnnocxk3T5S+PTMwpcisoApWAgaM7EiXsvyLRDws49Jh/AYJnN54hF0p6BYhc0v
enNjz4xqrJ8buqVI6dltJ3EhNr6TPm8E8I309WLsZ8rQTYydlE3jNWQtSHKfWJnc
/jWt4x9dOspb6FKn5u1I5tU8YpS+fBpn/8yPghrr7QnxhLEJIiIHRp/bJdU/EeNW
5MJc0PUurMZHpngBMsMBUla6pdC/dXFtHaZ50NzDGM1+wDIV75MUdWCqemAMySpQ
DsDQQUBaMwTDlNOXFQQ9qmi8Qqyh1uTo5X6Ol9lT8qyA96aggputcrpWPkoFEiDp
96MmAccKKojipJTVbv1XQ8OZx1AkgEwMCyeCvTVnylrRaRTb9R9EKrEuTh/ySw0a
K9MkyZU5BUFS9E0ohl5Km90OZ1Vt8tYc3VvJ9neheCYbwdZJAcJfYiPJyBSInlu7
KJBSJEi828lrxYX8obOzt+EoGJvDj9ZrtcNeDjgKjlgc4g4jpsL27hclT3vbVyud
JVTqTu1/Orel/SXq1uUoThN3egvclbMRyO3R28kkGLr/s2SqqeO9/5hC0+xt6rAu
p2oXao10lVh1wfWyaVh7nrUk1ChG3wxC9RNB615sdJTVfEgU0HffxQ9B2V4oVCCL
Q+qc7WNWWjHJsnDfQWklLLhhtffxPfTVNaDNwx5r8VewOYEC+T9i1GvQ+t+5u4Eu
bUZvZeCbooI5grDFXA+DSsFpNPMJuTVsk37zharks80kg72yguUAcrhslwBwQ+UU
F7ac1c7DZsIwgpuRwc63akz0Y1N3ulQyRWNYnLkerygkizr/ux8WBIl/7eE2Wwbq
VuUfqoZBgDgzUTUN9xpZZBlzbqqt9I0UtqTkDMjLrLPl9rdNzKEbAon21qbycrNz
cYgLm07yzyEPEp7ru3K7I8Dun6TkIzt2LxOOnDx/CQiu1zx6WA1IPNLvFyS45sBr
qziy8LDlqAhsxL3cax6Vv/OVZGm+ju/Iho7bGlotHPOlSk+aepVCFhCADs90B0xM
L3WdjbLG2aWEDjCBbrPe0FlkD7wstE7H0lj05bJeHJgIWwBhIGod9PCz9Orb2lfl
bYJvb2RmhjLDFRf7aoAMNITb0hRpEpwlvRiloJVC8PbpQkbPjxZkYsKQGJ/ieaAt
5ELq5qYrNr5TLl2G33ph+8h8OeceL59suy//SbMaWh8TZYU2gmrjde6gKLbtbo8I
XW6INxV+5jOifH3FN7kYNedqGI8Ilc2ugYrJ3u6Ekxcb1Zi41UXv/GtVLLYprlx8
ftmNb8E1lM+K+bXwHdfLTIwEdwkLaAigKpo8bdo7AVpG9wnA8eh6SeixiMCiXlKi
MZVl4UDWX4u2m13qgJx53pKQrqKYk8HqrGguri0awHqK9K/bM4k5p7GO48R5UHvS
DMk2FlIWvETIF6FQevgy9/dyT7DyKpk4rstXtuXcvgGY6B23XqK6DZMyEuPQQ8RO
2oBwEBR4gVq4J1rgE0px2KFT05YixagMCRwYNzwsqw1bNDTAMJAakkBxedZ8nJS6
I/AFF4WifjHJZL/7VqRehIsNHk8t+WoS0ydHZ/f1HYuevYthJWMSHfE7g7YNyOXX
s5s9DAVK54TudikbJIfIoX5tuqaZCeH/kHe/VSZ6/10d7tENHEexJlPNiCNIfzWP
Equ4+WOjlHVp+URiN+oxJjsZIEaY0iG1r8hbX42DJDfNeFa2bJuqpW/5fJ/nofBh
jWUF4rJmaTqoMwueUKl7ZEVadrBIE8Nj6vnhr5m6UbKXeFnJ18yTLqt22x9m71LS
WFQFnzF0soOYB+jGEJcGkPBUjhwIscmwNluTla/8XJoXkIqI7YqavIushwIVYwap
1AL8rKV3ChDrrDn4sCzGpyCYwNvfex+yYmSgxnKmcnfUnSL/rBql9aqvzpkrvu1t
X8/Fm8uKgJp2sPv9wSRb+YZALLxANH9z0xfSsoowLxcbLjqJF5tuEB680wHJ77/v
sz/rmIL88xq4Fy+Q3RJyZ7iZNf9MTFwF0pJlRMln+sc6LENhpNdDybuTOmY11WQX
uWP8ADCK0ymSk7WLZY74cewNkCYRWQPZ4V1v/yIQfpYKOf2yC7VxQlI+hpzxuzxe
Cyx6+A8HW/Ko7MGa8YwbUMo47IxEfgJdTEWSGiuWd6ySYVlI5ZW8dv3fqy2EDFNm
qa8UYJ4udYfkHq21LKMI3uycmT0NUlvA81RIee5Y2bUYo91U8kBbhbi35/Ohrcq1
oeIN5hcBjMxMlR2/CDYqoLpsJ3pDijtSoL2uIx2P0+pQ5m5IFMktA1GSmJGmU9cJ
gzNP8Xs/xG7lNMHGos2jGnVlh/5kprZzOHJAGOeu79AtI2X6kXw8LODq4ZYaG/Oa
8yULx7FwzbP+6pPnsGfR0B5FxY6fAnHgAwKkTvGDxAGOzO3E7nFTju381eL6K+cc
r64uhkDFTIQenYWa0gpry4xKme7HEYbYP8w01aP5bQlCO085MBkNlagWfbrAh3Dn
+cc1T29w8uSPRhkLiMQpWkh89RQNwcS4Y2wNig47SOG5+L5TukrW6/u4ai8hBTy9
ddHjCNGmoeyCFthuAwRa/g40vPjMZzbYAk6fqGA62p6YRzolfhxtJq866J3/se9m
3xLWorjo+P/i3Qgq/Ep2FQpLS49pbJ0SD9VNEc4H9RMqu81uq1Y6YZC47jpV20XE
qjI1m3hUZpSa3/gmvOQrpN55JsdhMTPixKwBRwNzzQk34LwGeiSC9P/r1SwxA2re
ajHV6nFqd+O27S5PswgIKH3/iTLd1EKXgrAPriwQUbz6sPIIRYHKvCciSfEebL82
fEK3+B8t3A6N7fNRgAKciXbFBqMfZdJGupaqCjfv0eEmZPUjsGnrECEVymsr8dDJ
xKFHbHwoC0hi9hkPK/dNgLTmZwFdM0q006d0hMKGxiICSN31rX8SVsaf3XntQBsq
JrWPyLtChH1FuEJw2jU/vccVBN77qdj2Jx5iiCVL3kFpkGanECJnXdZdkFvPUlW1
6nxJq6MMN6A/PLsXVMSmtJSq/by8TfqVH2NnrC44q8Uc/YH6veYyklsPo0bEg1TH
FjW5FbtLJlYTzQQAnnj8ijxPKWunehY0gs0tPkYSssi8jIhNETctcvbxNh3wHcrD
VLAWhp0efi6rdEl8wt0h3MvxuZoKnetKMlUOJfq7BGyLAsTYE//QUcU3gpT0Uovn
SlsrczoHbMYYeiImDWrTqZhogAtrBVziFAz0eLyjyrr1LUbgyDznpmmSDJEXuQS7
M9KJ2Qe392xR3bHGTokOpScodIhSyC+IYEW4NXJFJwvTAf9QvySIu6vUgJYylFAX
neguwwqMyAsLwKHYW4xyCj1G17xfMbY80R+d/HN4FntQeK2SodIgYffzsbKVz1o3
hCWJaM86z7dRmLxdnPpz6zAT/H3FFW5ZLEBY4J+JvXGcFf/6u+GAyvqZOquMsJeF
Ca0gZVwlWf8nr2T7f8VkUw6Ioj+q9lyhAmXTwYJSlyhqBQLnrzwuKMchAastsR+i
tUzr4JciANJikbNGEv4eEcNHu37A5Qvq50AfAu+QSFeUwSyyo64tJLv1FjAP42Yz
2GwDYOqz8kpEuFszMmyVm+RmvmX12L9vCyaYzOUMhnXcAVKbj2fOKMneZ//1i6at
2u0QEJT08lMOs+jo6h3OIXmJrXUejmKfgN3OAE19a+BsqV3dFL1fJSQN4l6luZ7X
1yhGAAp10+GS8v16rxaJiQGRfV/ghDapg/xupxFD8AuCInacSpn63xfXmS1UmRZo
3Wb2glYlk81TS2iAWyuvQ2Dkneg7S4BPgHYxuj4IqazGx34t9p04gutodjFBZ1FQ
tOZdVyPptIa9jDFSqmUqtZVUc3qwkoDAOP7F+TYaAMIss3ehwRtDP4dA113EJirn
AEmPRlbz8mbwDJJ4hC56EOKVdSpYTKqktdz6WDdUCZZ1tPoAf9Wo81Xn3ZTrP7Ir
nVtPXSCkehq/HcFZbzvj57MsY17L39NGNzOsW3KowGxj5IEqt2UayPufzD9j/v0h
pqHUyv55wIwyslaNeNGWgG5yOSdWQaemKXUPmLgMhhpRhICpzmvZVu3cawLvO525
NQyE8rSZ5yZBSlPk/cZsIz7MIY1oCjjXIexGNHXbHnzwZxvaPSCTQwKJO9FCJCb9
loMs5G5oR2e8Hd/sqLTjK5UD7j46RQ66L6Skb6JH+Z2vvtUirBp3p59T40bRU7G9
K05wT8XfhZ+OXhxlTNuAoFm5nDQ3jYq+d+tg3BYDqv2U54ihdraV/bwev0UPC1MF
wMI/y8PmZG5R580ZADMcoCKubSgBdFkWbo97Gk7//tkGio4zX4udzm0OLt9VlBx7
M0Ga5Ujn5ATzUTNMQa4MTC1/PEloa58Wwy5WJeM7n4emrOrAq1qFsunVg8HMfRVt
kE5dq9kyrTcXY4qf96uiLgToNX6pH+6Ktj7BmXVf15N8eWjIySRqeakh61lT4pQO
FMvuuQS8hxuZWunILVGZBDAbVqoVAPh1YyJHkvADUfc04k8mldQsFWi5PmK/R4eO
yesoip6DTY1umNlBONfb6uij/LEpONsNVf4FREiuf5dUu2qV93mR+apFkJHBGviL
Xuet/stcHtERISbWbIu9HS6jU2glg49ryOJLpSjmy+MWtcRiixG6orRQ6/GMEKEU
9IE0RM9VNVDrkq3HCQM+Faf27lXzw7um3hJS1NHrMnHX24/rUv0J0YR+NSEK1dA/
242gHRXj0FGd7VQC/cq4t6VueBO8Q1CqlkGd+YFHRL0xLLQ+Rr9UGQvHIWJz5MRQ
hgSwqr18T3KvGz4Z9YHlRTY9xTid/Tvf6LiCBV7X69l1v5qPnAPAkcrB2BnzAVNh
XRqnHXXdnRjyqEN12v2r2mMaH2LK4FVb1pRfwQ4Ld24DSz3lY48vGDimtI6iISMs
Te9AdkYOVzHcf/u2KN+F0c6fFJnMkPkJhlkJSHFFv7l/xegmZh6T2tarTfl+lzlL
6R/E9sqDlMR6bwE4yydCH0NOWM973Y6aIFg+OxlIJUWhmu1EVD4fS0eNvTK3aJQ7
IGVWnXIJe/o3tkCcVuE3C/Ma/4dHfpxZvSzlq+b67AzXP/hMJQ74abqO8XYRjWz5
s6K+XBqybLG9CKV+oYuq3WP9EyODA44SO/Cn/HUPys7uUdyq/AiJwUVTFVV9nert
tWqMzWurPrZxAx1n2UGm+hj/S8uCGPLlqVVilHrXsAgixkViT0kBFpu+CWrj418F
ktZCgF/SmEBr1izPlh0D1rVqvU/0V0VANpomUbmD7TZYJdxJwldABXqaLN8zKCbx
zaWv3zt5VTwj5p20nnC1qQbPLfPdPE6ymklD4ovjMkuIR0jUBy3lqD06G6VqCoRL
76RLZ3SsCHvmHK3aagAuPDb8bKj4x1A329cEEck1nbKvdaoHA6L+MA5BNd7/cFTr
AoBuottQw+4/hG+lvuhlkUubCLXwHIF2azpaXQS93i81vYcSEqrVPYud+RHG8M42
taaRXIXVr4CDLDGuHR/zbWn7kzM6/FhyEDOsFNFA/veF+Dliu0CGLa70RosmcYri
DhYZ7azwRkWuPE92TvCEaqPZvH1BnnRuzTjSBJpiQzU3ipnbI8DhGhmCXCs6Wrfj
QExzW5HytPmMRSaLS0a9X67xPfpZ7E/KfW1a0mm27iaEAv2rcqM24dVWg+wu2Xq9
lMEmXnwzTXl9VdVI+ow4jaAd4V4pzu3tvKl2HjUdCBh2x7CdmV9K0+RIz74DEKbC
QOaA5gCp3+DEMFNL9/jlN5GDKAG9AZ1Zu5G/v4WrOz4wozuIvxVvEQ2j2dmm1qk5
g4jvGwm9izA39uSQn/iQ5g2Jve4gMGt8QtG3wzYT31ZukNyPy5ecu0ta5eg0fj51
k+KvfbqLyBtf+nQY/nF6DFNoHIsD/MRB6SNWowG9bsM/aFtKIgYlmQox/KuJDVym
6rvX0Bt04ZMIbEXlJZL0zqqVx4fNJofbpkwxENZpaxGfxH6qhiQvLaS0wwuQBe5Q
qRT5qSMsjKGQjmCP3JvphfLoc8lv+KT88UGT2dYMz9SwqVfRMlt75axYBFDyB7QZ
1tAeX4RVf8o+6CNgHHmQFGWG4jC7JAX+np0I5YtjfBtkl+Sh/mZ4ZB4v7Z00Tvpz
+1/WSZl8ErbepicS3LUlpKPFDcIyRISpQpGVzsc0QSRw0Scd8nFw2gbSmYOI46Et
Rklx/e4UrF5vruwN+YrZGs/7xSN7a/OfUlnjhaAyFcnNa5IPrh9z6CWuHlD5Tu4e
B1mR54D/Yd2geKZ7dOCRTinZfTIKCG56JSYIKXP4PA8uvq5rWO+Qw6QMzLhfdPBu
Aiizov1mxfHIm8CEHGu/9Im6e7qSM8d5zvDdmeB3DMwOdPjhEZb/of9f6yDcCsQx
Zy1++T6Kqcm3gGR+6iGmLNmt+JhWDWTR4f/j4GE59FeLi+mI9YPFU/pBVAprJBzw
DguZdzXxQU8sFhynzy5Ep03yObvC9QAtqxOrGkopBycFx076Pqyqeh6D24aZwi56
lpIw2FQqy0R7+qLxCPdMNrZGda9RZ3YRoYPtkIqksV7GqMMFocddkzTVzRmCpr3W
VC+XNv+VJrzPAaa0lufdy6b815YxRjGD5YCrwdORqyYuVobWd4yxUiYxAW1wMEtz
W4LEjgd+68OZ7AcRSv7tuERhBe/bQTvrUTom63K3Val2ShuWmoXkrGSy8yZnYNbd
nEeoasgA7tbo8HScKRROS++3BafdL97wCPMByy6ul00qoERqLl+hNvd/D2YtF62K
fUw3ZkX5M3lu/mX08u+cMcu8frsSt0XpJKb8Ziulono2LPlLE8kZ/Nb4CdRZDhDU
iYBCClUDkU7HqolB0rZ6TSK1a5L5AmzKY8nTXpv6fbl9e8TyZjDlt18bBph7WXeH
7m8yFC4gzVk8up4Wgcj5poCGcqTVhWjPTMJOE5+b36kbziICBIJx2Sp/jqytkEJn
JVQFxcdAzlhXPqWaMp0edqz992m2Pp0OI+rm6eiOwu195Ox1Aeb9X2jrxErOMgv4
RTo1X2OqaPWTBwfUcbYxdyqn8rHgkx9a3++LGpsP2oZ0nFDlXUfL3SPXm6ajdclV
Ybc6sL7m9tvxad+9ttOGVJ5qXmJV8G6KfdnkG6EKLNkmL9Gc+hhpKBgSb6VVeMrO
+7AZAe1sEulTkyQOcG4vXQiOJQ26eYrV412RpqR/5fnbBeqIeDVIKgL7ngf+5Ah0
pjA1bcxFHCNfMYhvA9vsoSOfzzoC9tgtbV96XKUIh+mX54tHGsDoO09/5IZjnjMC
tm9BT3PjHQa8hFT3XHoHh+ML7XG2fSsCzydpcnE9DkDsb6Re6NwAKuw9/IrabEYa
K0NzLUp4z3Tl9cxg4OJJBlncjfZcqgOye0DCfzNQ+vq4XiZ+k33AQGuO0JsAkeit
lxW6ZOAIFOv1dB8Yn0NIYcbYlOObjhkVUk6fgS6KREDrWFCxmhX2au2jc6x5byK/
X6glBHl+DbqIIBU8KKl/2NeokcmcsoiZwYC2CNa544+HJ/e3t7UKE4i03Vcx1s0T
anlV/FSoaN0OccWHDSYoDVaEboP+BnM0jJxSVzbHgMY/Pu1BEurmPyG7RtNOYTr6
i83NgQFcLn9+0hOvOaJUuPB2D/oBpPCZmzX8wyawWFtMl0ON2yrBLz45lyc//uJW
darISqM+kvE+zbQ9DSeiIV3+0WuSfAPmVkm9Drp1FsjMU5GEyLTKlH3nyZeVsXuB
8TZSOyCgtgBagHgqP+7EWgFL4ImBoMmsgl2icGE8LKVWYRpn+XsAiwkhIkPFBTNN
cy+WxCP8S9os067O7llJ7MdskIel7pIme5NDgwXnsbcfgHI45sBZPtW5cUMH1HxW
7ARr3Js1pExk3T8o52ctgnES9SkgbOJ42nuGcJMICNw04RbOoqWzBUAZ04Typ7e4
8pZs8hyaLo3eRB1/nOlqvDRCsZzoXoFFx2y2MS+IvhXfYJYPmYn0D3S05vplQ6J+
bE8jygHNQvptazYkFHJOvAvSy4dcmFMS3Iy3NR2wShfEROUBXDYpFgNLZybKcAtN
VNKuczSjPZwVDPicDWtwEw6rVmU2QNrA38nw6JXJaLXrjzy5zp7bvCryv7c+SjNU
yJ28yCvMc7Q/wFRqVzpIrLwJdlejgTa056H0tPQJGrwoIOdC8K1jGMYAQ41B/VTH
kZETe4OkCja3ijDz1xtlCajklEvZaHaxfLIJX1z5s61UG+IjTDHnZFvL9M9L3Qpu
We9lWpt2VnnSCIVQcH6e8N3Upp4GqJhn8oCRKfVAVNR+KE96Vk+g0+IRFywmDdMu
dCpBqq8LIYSKzIz6KnJ0ScZHH7bVY2Rlz8pGhkSk510FSh2dx7YTv29fu5CR8nA6
vwYlN/ZwQAK3YldTVzIcfwia23YmrH89SBOItc6GUwgbJMD54DZ2TGio+KiQ/Qd0
1mQIfTs7+c2UDeA7K20cXC6CEt1hHmZgKZp4ID2xp45E8ys9PI51GJ5U4mF+Iz0p
lVq6YE8FXgVaw5gy9a3OFRtZZ7y/4Jq4P4T8jU3ZTZR7H2kHsXexCR1iuNq/0JOD
NveTTlw0WbjJIwkAJ3+v7X9dU7srcfFyuc5ITKFyNkncli48L+XPWB+nTVKHdvKG
w//P+/6DRdNuYoA3aNvu6DCQjG8vl3FoL0AJGODnkyDFTvFENify5d+T7Fsi8Epb
A4Tk805TXMDNs5Cn4G4iyC6MOKImJj5QQTIeBA1rndrg5jcUqt1RtZPNc/oMMwEc
F1f6fieD6oqQLFNKxvjgynekdXo3jPgGkai6Y8UyUZAL4rLIo4sV++AET/GWjbE+
3J/3Uvi4ISfbp1+CmqB9b4WehjMcZjpn48tSUGLbWD3QmGQB10GKPJEv6Iur4XKk
jDNZJGp3RxR5I3HtZpaRYnwB8/rldyNx1c8tpHDIA8FoGAgHEJ1xQwp2nzvekc2z
uibg2EyoD+yjLuo5N27ejj8iyhGCS5eyTtMdcCFyDqNo7lw6zDN+iYvQh0W3Y9AJ
+8qDvt/8XUwqIQMBBWNNKgZ3+l51rT04kD7h3WxtnwsM2DnbOZpsXxeMNZjeZogz
oU5QAgvqxD2MN0urBRaQZkimVCLIRG8X2VRhiW1v6ZGdjUJQC+LmZ1qnN2FjwEed
G19yN68K3tll6aiHKTDsKR759FLjh3NeqbHmXMDuyzZKR24pLKzoX8sPnaFSmMAE
n5Ri0EVXWfjyCrjWI0tkzN2fnPOmi7FFKgogUmQJ5Wsm/dG8IIOPgOZz7Exq89tO
6Bb414f28PEat6eOaF1yIn5NaMFX6EeEAQlOgwKGfEfxbD84qlXmyIOuOPE61FQQ
1TgVGvzumTMz+6R1Bvjlod7p1KP9NmzbXAJ+HeE0HacJU0mK9GM61fNdNJKSJgJd
RHRS8b+Pdts2K+8LlojOli8Y2JGm82Kjjgp1GJngDyDzE8Iq958IC4hv1IKoK9gS
0elYkxDfsC+abE1W6hvf6sl7khxONYr35qYWbQzfsEPcyztN5t+ZwL3tGXrhRNnT
XxCR+W7BWgyqTSWAIwCU+VnpSKaBqIlsapXWi/BVrCN9pn076yoxXMTFK1dt8SWm
5QlrXUIHW+G8Y5fx6nYy0zHFva62oIvqO3FyKA+76AMCH0fW6Ihun+23yoH5Aaa1
Qtg+n/mKPdY8rkjuyTWJzQkZf9HRcWzKJgBa2wjlXg86TYG2Fi7jMfjrWByzK4LL
T5O8eJFlT3XA+kcWxtfxTElXFuJAKdXGR2q5aAZL/qDDSfF+hxqGPGb01omtsfbJ
CGvR2XDvw0ooItdI6tQAjG28ZZYcqsOUewl1hOros2r2xQRSNKDX3OMpFUMcYf3j
nmpu4dz7zvw1zm0pFmN+iwQ3S/hnvlt1+QSkJchJa/SqGtxDN2C5+bYi5N92Z1sz
KfxcCBOX2omUOjCNlV4lzGfHgYkv+x9TUJIAXdW2ey8qjzlp5EZtLNnLAhCSG5X5
X21HVGyGZXLpyd0hSYj+9FpFOfjS8LJ+dbEpTKEVn1fAdz2F3b6zz+IX4m/6B2r7
It6yttHJDWGBh4UFiXyc+muFWPLD4CKuqG/RKHQY2clSuUGuFHTX8b7tEndt0gQC
U8p8dKV2gi7KhbEfIvPYZ/G80jGqwcIF1mY2IdcFkCYtOkS8lWVMyKDOUzYBAHqx
xL/p7lP5L4dc53DJ5hwJgV5a0JoLotpKnAzkRZR/MA6JaHEX4otOCgBxYL/DU1yr
iR9nUdFiywPyDalDBHGHkGicW2miICsYie5Pn3ZAKCb5Vs8GUdt4KNGeAeWY7brM
erhXoTB4g0LLilswj7f1jF27j11C2opjL2AUx19+nx3MRtTsv/w81Kxnqbyqn4Pi
GxuF5BSyBOTn+miVq5mwL5NR2k+UYqCeu3HuNwNeSHVvK381JlQ0W3pCa2O0S7Co
fkxxpMuMLrF417u5ugKesX/GHrdsr3fo1aYlQeYAKOO/99bIO0LoGm8A07robuHm
nYFlI8J6dFyBGQ5zHyaEsL0nA3WCCE/98u2JXa6wyxPAgOXZts5zztr2kDcruxsV
hZOqPKcUCF2DEuNR0pb3sVFtRglj8fVckuCIYVz8RLWVYgxgy2uHiDanUz8TQJEZ
fNUIhVRrFXX9V458oDoeKlyOGrmKiz7zuJjKzYRCo5IwdCTUiZyzthvo+nvYrwIv
V89wbXW1gq/ogA4qGAD5XrM6XAJ6aRmq4/I/mUmDanxzWoIZTr1xuMMAxkhIlWBM
dWgtsNti3+HlDpI1zuET1BV9gUqg01kkA2EYGMxOIBe3h+KAQmF3jddfhg/Rqauw
A+JrB4GTuge6WjztVR3xdhX5om+5lzoUFvJ692oxhnT1+mEbDZuQYvfMBPx2aMt3
XKQQQfcE6Ad/GehKN1xdlOcQn/6kUO6Rwcspcyz0k68kNnWn2msz2dTjxX1SWNYT
5QuVp+HJlVq8SwM2lPzJyLaVQgfw8tjKW4OGH0VEdNWcKghn8y9cDNU2JIu0QyGY
ALv8rAYDJ5+twXBZg+jrRAQm7l+z8LGWsuny/HMtxSxouR6rM54y/SvjYLUTNtVT
tE1EVpW2RFGBHi1OI3pOcD9iu9+Wy2OHgSFW9wvNsdOHraaj7KrZzhzINnvrDIp4
a3Wf8N08kTv8ihpu30eC+h9DdlgJTR4q6cpc8oBLcQ6vHH250YcsPMOFPpSpm5N6
IpqcCxuf1v1u5ZFkbm/umKGpshwwIo3UY7STtVlGdAtEONwbsvO8p3df8dZVOhps
rBsiYvQvoSKnFM03XY/1ybN7j+Ql+VSCbCr30WS9waiDtRMdrvLyCNS0I8Y8yVM4
DmBjxYJg+E60SuhBZgv0btseHaccnV7PMkrTrH5OYz2FotLNkwGv5VeYL65IgLvk
ilXf+7PwHlBMb4WV27YFeNRKj/Q4dHbv1KT7XXJGCKOZjqC8JprXsWLy5Hn6k4Ia
2Gs84TQvq7ff4lCRgySx40v7GDlELPCGvevwbhNlq8AmWddrLRo+1/Qdkr2fSA/i
F6ekGtATRinW0Ri71EUH5V4g9ZjxQ934O+pEfFSJIpS6RBkFkBQ5mpUPheaneqtP
rb1IcjrAK9dlwSSxatEt40xSriQ+zsJAJqnzF5if0/eIy3dg+tgJwKNcRqsFEbHc
1adjXwN0mP/DLAbe5v35KpCusja/QLYyMQ9g22XmI0p7PlfbVfrhvA8OLJ8TgWV/
gM3g8DpmOVTkQEdnT1nScO/BJ9O/9K/xF+Tv/P2dr8KAlW2kO5g+F+bs25u+5wcb
6XtwiFJdCe4ryfj1agyAIeQAgbsaNSWZC2CjYwyA55droPwZKDXKKOoVcXGgPTP8
1j0di1Ab7hmbBoFJSlgA/k0418J0Wjvr+C7DkpIFi5PrEgGBLTbBhwKM88fIxTl6
rUAN+SX8TyajlrfewHbV50wvAv1heY8aGb05+kN2CVL13/NX9UKyuzi8YfkuyTa+
yQScsvi8hteBZ6sO27lnv9nUy9qm2+60YUT7RgJOx/zQ3QYnCy9nR8Oh4TYz21/O
RRHERwNbS8PUQ7ajILk9HWAskY8NfMhUca5kkBjBGfMaIyRwTPI+fEhGxnXw0Xup
DzQrerxaljkTKGPf30Z8hyRo8GPBoubXLo8AHvXB/HZeMSFxp8tKI+ymS14wj3vi
KBpEnpuFcmh0RD+RaWlN3akZNhkMOncUMg84sOncZpiBupnUhr4h5hpUM2bazo3p
YxDd4PiB1zP8hgxkPOjB8GSC9f9SOyMCqv2VCPGdyX1DcRCGXjMW4pMI1+01aVH/
HjRYDJ3I3WMHlbjR2u8ZKAwuibTO4f0OfJGxdF5uZYS53IPuDdBMNMureP2wzxw9
d0Dm821krFIzpc+bYX3O37sFierpA+8pj+MK2W/F2zUd+WD3St1VKOESRgeVI9eb
fORl9BAgcT5BLg829tDT+obEHjOYUo+ZYXJ24ht3RZBfoO2qUGHR89HSWz8Ad+uk
hUBqCf5N/8cSM4QE4KZ3i0DCD1Cp0mPS5PTSWE26SxeQ2mH53xJ4Q6qS6y/HZ7lU
u0IkareY4hKCObCvMiQcXysdbQDa2AjKVG3PI1Y8sl98J6IS8+BRF4tJpN+LF8pj
d9+4AuKyWIDxyBRxPCJfEfkaAuxwGtw/anrI5eNZkLJr9RdzkzBytMb4wvQoGWd0
5ZdJqvFDOTZpYyK1j1+dmmA4LkG2xanlkWS/wy+4HOsL0TFzfLJq4hNoJR1HNV4G
4OYBkoN0rlj5p/LBIyhwEM89vQCAQ5QBOUxUENolezTVASidsghtEpc1K0Y6Z2JG
Poe9rTY3wsfLRtWAcdAAVlKKEcknfDFsIb0TfdOOT20PndRqdbCMtwQ925Ec+EGZ
YGybwPNud5gPpiOt+EJoZm1XrW/2D0BZZmbILrdW3J10N4641UUE4ciDR8aUyQH7
nPC/n5SF70G4Kv0wyDKYssoCcV7My0IAoJ6Wsuz4pGYqYg+mBdoZuQ+A7y+sVpfO
W4818H8UTLgFJ/fwoK6WuY8j8Q2HyMPr5goIX6k8fZUmfaNdLGVipNknZ/rntDUV
GzUjHjYUlikj7O3QkWvCDDcgVNU1K0QuFxCPbp6eLpkD4a5m8fSHkKTtf02BKLJG
fm1hNfdYvjnZJP6Iu1EYjUXtM90UGXlzPEbuPkg34m4uCRAYNCUIU7TrMHLVGCMU
fwiWYIWMqvLacO4J9ii1PeTrSc6oo2I6lcbWGLyXWc6NPbgz7qAPtUSidGBismeJ
C8Ck8s182qTn5cuWRuxuIevNNuDO+DtyBohiW6PgRqEHNaeDHUQ+Lfm9hrgWgqSk
Iz9OzZjOrfvWscy2RGpGDK/Uehud96+TA0WDbS5twL5Lpw7UwNskq0B4HDJaJOSC
wUAhVxI3s4jPAVxZFn1y1NXXJR0XBtYsN0IQRReARhIlo4xyn+7LFrasIUndDVlm
VH+nWlesqXzT+NDKIdPLQyWz84vwaFfe46xI/Fv4qJiM6AaPgqKGuqC1SSxNlHmx
vREk7X/35Dd/ROimBrJQUhEUte48r7u7cfXom3j6szGZ5jDhAIgDYP+OMKAQiLmA
dx3yISDpLnlWCvGraQC3cftiaaaQ7ez1zDJ9oEiQZJXRRAOGbMPexQiKBPp3Vhqw
PY6ngJQ4DhKejZmyX3+G307V3T6OVEhafSknrqxFaMIjdp0LDNC7yhXykEekNzKW
IiNCVgar0eOx9ii4fGj99ane6hNhWeOJHHYu1l1qGyczOLVsQETr/1z8A4V+SDIq
e2I/d1CP2KKPQ3XKyeZp3VVrSWAkSpAJOzQnjqwfkrjatJwar/x2t1jHaRKXgusb
ZC2gYihjf3veH/smJqI6DQ3wyqKCdHchSIXSbmE69rZKyTQWYJTRIhEH6K38ifaW
zACFDaOsSk9E+tDUUvTW8nQgo5W9yZpw3ZimcYIS6GdK4plFmupKbuRxJJVIgFVY
ypZ2T9JJ9DisVZBaf/5ofrjYF0gy9R1kALcfW30ga2ZHuyZjLlrB+X2ePjyY9bwF
YXAg50E20QY62aEgzWoTE0cCRh6HAXaPSzNsNEfKFctYh4lattGkV2KhkfFz3HOK
YUwQrHABrgbl1B23ERezpA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Nk4IyQvuNRE2Le1IGqKZh/ouVs7LID7ml53+HJhA3Q0wRvRfRP/IIOwmNZchPAN1
WItGx1g7gvp3k5k8vxswZw8MvQZCnhKUOLTp/NekdWBAIwwFCf22n3HNVubrjawf
orEW1oMUqwUPPSD7UGuGjlewprglIKOYc4ToyiB0d9HKcqvV5c+BZvmVSEk4vzjm
AJ9QrwmcRhz3MMCUOK3gI7+K/p4N77Vteoelcqc8iS2vyZYzj3oAgdL3N2X+Wo+o
MmPKw8blK+oOs9i+MsxMpTRBgtowLgzG0E9Gguf7BSEKjkA53EQt89i/cKi8kihO
hkitL9V8Mk9TML4/A0ErGg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22704 )
`pragma protect data_block
wwJPrqXsOdwzzCP9AxSnv7vODJCbzWNx2M//jJIlITnSRmknlHWHAPMwG8OXpift
zDz56CYGFddbdNiwvjGgXCjZbSSrpgkyBvwdMjDo8MrV+QY8+XlE9yIY8T1GGCyo
d9XyMn2RX0gkOWFDafQoEFnCmFgQtMRD2ihaB1zuWvdnsLGKQk7OVV5/2W7BmKKV
0jOTD/TQYI4XU8g62/jEmBFo+8gHF4gVapHrhgt+b6iNJdP5np1fyL/dKCgFazwR
26YlYT+eusmJ2Bjyr+w7eVanjFsTaSHU0qtmgAlovD6SYWF1sUHpVJjJxL6OBEC9
uk1bjrke/An4qXE1tRGKgbBsZkKb6MJ+DqnwjysxujjtbVNCIzaCLEFPxVrAuUc0
mdHYNhf3KM2VhVZO2Zdob51EX/izynbYQzVibuqa2JO8KGb+5MlsGGu/ggJpCHHJ
6zJXdk9bglUkjTlqIDN2u1M1/X7UuRBiY59s0x3vlAxL9uFlKz6DdgHyls0+aX3T
itF1zXxa1dGQqdtfGVxcBNdnF+ubov5ODJcS/fRJCHvYVK5m4uLojMoc64wCzSPo
nPWJ6GwCohlAw3SabgEKjYLprx1deraXXJeYt3DGp40dGnvja3jy0fWyT2NnNO0l
RZs0S/MIZgLnr2cYEzGCUmEWVpiysx/d4GuCrMmM94UgnOEtdzxpO1MwsYRmg5qL
AGtRDEYsXHNLs0yc1lSO2+spDrKD1/G2ojYZyDcv3gvlKDkv9cn4FgWGd9/6xTpH
WMyXPp64Fc9bWDjR5lxb9Iy/2j76xFuuhZQrHo74FxmY124S3T26dHLE9HzjAN8P
M3M7CI8PeKxma6aa8WT6vY3gRTAJ7+mR2L/2LG9elvCUAsNHZClibxSnzonAA1oE
cfcCin4RAUsYi+lp4eOcZuWEPwDX2kppv6sn4lW2n49k27Q8vQyJ37VYfEBQXmPe
2jaEj9Cq6YVINlJuooxUAP+OAgvtcFe5Kh7c2iv8i3m/3qWDW+g41F46CAoLSJ0G
5VU0TgOwWAkX/wubWISbSiPPO0yzvV8s3qJ00mToQzMjWWpT98YNt9E/eHhIBLYV
ynn3TcpywpNN+ckgJ7XQtPN0HMY/uqjh47mStrc5MCFJkJZSTiUMsHc0V357g4Xw
ZleIsPjTrgHfIlwZfdpLfbJcS0L6ui8ihoEtopv4KKv17HzMZlbZ0i1AV0yfWztx
Fsh2oD1qmscvZUdUcHN3cvkcY4yzGgCzZUg4X1eLDOXuCwbOQlZeYTW0BVk5fToU
JQKxG7I5Wtl548IFSihds+E7+t5BA2cF4ynVo+kHNuk6aKreBRwAl5p7ZuatyhiY
yA9cQyV1WXUZrj6707o0ujyXrmfoH8RVQY+WX0tlmK1mFxTkxNWwhixDNQtJtEAx
/tItpNaYyVm+IJzgv03+7PEFTfBjH+JRFjvY73bf/RNn0q1IuUkmGXDs4uhwLiJI
wujJxegEh6KJq1ntJgNRQH5beiQRx7/kiW10WNXueEexeN8NNdonupHu0ugW5WQF
p+6mbpvyL0uHkiC1OliFus4PptbDxLm/H380/Z4R5ns4gyPF3oMGf3SJ3I4nN0Ah
uy3HAB7EiVjDlFD4eQNpugE+wKHJ9FfMxyiFdHBr6zAyix+cnDbo0Eblxep1xtqD
vwbYoYRtIwjqMA/aUtXga9HWEh4gjBwI2LqX1KxMX1WPonr8XhEGP7kciVV/PFc0
XJ81WxKQ3lkod/h44AW3VPfhG5t1CcqZ/D+Lo4qDzjqjsWhL2tU1xBj8l4hz/5Jk
oKjCk+cdM1Q+AcVkorl9rtNJYkXLa8kO8rfgQKdr/ihXz8I9f+x9YeAJlzs54sxa
BFCV4XQ7FuDX4DfWpaYhdOfPv2mKubKK4d9MYpFDT9tAnVj+wpPdS2Ir1afiFgLD
bVjxiBSwYQG8CKQJG/uqC50U1wA6Gw4xI0lyNt0GsZoxqTgkxAghepnploqBhoVY
3RcrMEjQ/hhHc+gooZwQTdB2Bi0aVFYDSDbITwe3hpY3rlAu3KVMoFLKA8tA9jix
ySQlcqPuGW7DsYzEdTA5V+QrB4weapLe1KWi4WftN5D2B8fdbKobAROAPHlVQlkc
7U0bXtx7f5I5hx/SdGO5RV3utTxHiZ8x+1Vxz1mZLkp0r0qmPX3nn3LD2Bcb/gHh
VrnVHl4lSdq4Y3lr1kM+cA2/AxgQ353lYBgGWm3sD6iYjrUiwdjkm/rKZ9SuU0vw
htkff5CKqfYY76WdGoOQcZhZqiqbCTDbUUEOWdBKxdjc0qCmo52eoBsPIjSFaBrO
L0iBszN0Sr4WSyoCtLtoP/8otzcHjVheI3yXz7JIkCLUzbrOHBp8atDwj+GfA1Q/
NWlCU4+xE33Wja/YVpRaKD/miknA1WjTif9Zt8JpqXYk52ilAfXWCOAKK5bs9s9+
3DYx3RVBP9BBu6RXW/IBQH/nonxLBz+c7/kmvk8QIvr7SousSiC/BmA6Cy1hNbDx
iSLQMgLMTYD50/Ip+AqaJqrZ2qqigfykpG10rGXBvv7XM7p6hDjxwQgywaWxWqFp
UgyLQrrPk3JXKVsCh7dKOJ9KcL6AkVQgW0Xe3HCs6ac9kVjBfhSeZJ8eIBje+7A7
g6kxRaWBiUhS03Nl+pIwefRTDiGuAVsx+RTQDrNwEI3PbeRooHVP4zYb8tVfuabf
5f9M5T7mcenijkMADKLCF9PVMU4U0m+fn3pCQWGLECyASWqtGGB94E4WleUFMxKE
S+Pa6uF+U3maI9vf6AJ5BRedPxe72U/TP31Ma8Ak9h23ejeho0vDyylHd3RC9tgn
nAUByQ0KzTKoJB/JTz9l9cLnDInBeQ0fdSl5QWUIzIgNi8ALLTSikK5yZcun/2I4
adS8EwMdsz+cVucWyQ+cEB7Yg5Fnmrt/ZiQ+N9mB2wFy8rjqKYA1tpxD6sOtl6Yc
5xW9Mu70Xs8ZUvP3ZhHtRXKu95h4VvS8lOyo1PIP73TbG0Aw5+pPfR+SQF0fXnSd
ptYD4KTwRqh3qtQCYcGk3WgWhj9U6EqqWERZLP0ASrMikXqTkt4mFLOHM9r4RBaB
xZBeFlsYHeMPdHugKWpKDd7fxQBYe/zf5TcLb5zeui14CnpeBLDOr4VtXC1xyr3+
ufpWIau8e+150y00yPmBqr7fOxB2pkK0FWbzD46o6kSnl5F8I2U03L13x6avSUx2
W5PctIPfrjybL2Hl/K8xKrO68a5r6OXfD4KykdqDu9/Eb5scbNrJmfXQSkyGFAvu
gIA7jOEJ7KqxpR1C+RM2UNbKPy0JweF+3OhIEdtaWCpl2EuWv1xJHfZzmG7ZspQ6
yyYlGdwXEGh1CdjfsUGAl/ELfOSDMgnCnqMTvNZWWajr4ox7Eq4xHlSBaKqRd2H/
RZQPfs7oceBuTCsw5k3LYKEBa+wM9BE1P5fPeLpaNyksONf2AtQanowYkSbTgtk/
dnIAqU0wVEaJVAsyaOpspayq1vFASkqRG/Wb6Bwqqc/guHbDFyn1lsMLZputg8J4
pcDh3yh2dYcb8F8/WoX9fqzrmywHjxloqFF+NyPY8mxqDIxDnM6UfN94yqqm5VzH
40DuPuTn47bHjlv93YYG+WqSG4U+drxGvSbEd+nt01FURpb63MSMIkufugTuVjc3
GMek1RVYWpQa3KYQdIebMR9T37sVN6b/fj2YJbTtgOvHKsh2Fuybfdn1kkaw09B2
SiVsiwl98fQEfWpIEQn6lA2ID/oMGiFLEyKIzFzzmgQBvOpRZzwZc75cZD//wNJq
DPk2N9xvyyykk5OS7jwiisAOZkrYnZcxdtLvekPulVYC7aS2X+kG/r0kIR0wgK07
iNhdfAYgVI2LITl8F2gxmqW7CrUyk1x+Y6E2DE/ZiwUNI77Aaf1UUGrum4yxBGqT
nPWfml8kcKfGqeaWyTBenWD+zL8An3ri28PPTfyLrh+pgZ4egd0OrAJrbjxnOdvo
Li7hgi7H+2FfkB3q/1GnyZJmctBOFimSU+CFxrnppkKeEzf1LR3CsHrImlDN6Idk
EnpzPIEeze0QlwFBx59eV6v+67khPCHe5SKI4rM2Z1jOLHeRqSZzmkcNKWzwofWQ
IhwvLvaO7VrsZX1DoM0PH0M07Kmgc72ZGJif46GscLWqHRTgFFrD1D/v+F9xbV6+
i8VZ69f5n9L7vbe9F/pEWuQPgtf9rf6dzKNsFrltL+DBi/9ZkAjKeB61cwSw3KD2
BgRDr/456zwhFt01TS+TcBmbkObt//ZRczrYCIiLc0oRLOE11+i+jlhc6BoIQO2c
F2to7MHW6OHbJ1zatM1v2J+QCRlpookrPL2Npien4mAHJ7iS5t4h4OL7Cech3gnH
Tjyrd5GyplXHS5lDEaOuxUOkEhwNeXF7loEk2xkovH58CKgLrBtHFrwPR28LOBHF
C7b2ttzg5l6jIF78qgTxRAzBXQt1WxgpU+SK+611a3iy1vuRi/RyQcXImgRASA37
jTWPO/vm7pnhu492/z8P9KNFSLGZjt17aB8kL77noa9ZNbBqCOQcKyZRwYY3aXBf
iZdXgzssWvX7rRiCsWgkterB6uwjh6N5n3DQOVYUxCXxtRRW12ybs//tewcgqXdI
OQ6Nt+yJJFdmiFkQ1O1hBqm8ocW83jepQxnIhTVsqgJK9Ta58Otj502a7RYl8vOx
KX3tOAoDQwUN2LqdfjcUJGl/HP0fnznhhJY1/BGD63n9+OHPBx58rEBFUGehks/7
+a1vFIMR1E/mWNKK7kgXICAWjXH/6lQ26x1R4Rz20FjxKQtcG3Tk0etdcxPxu8TT
uw+yc3QWyBAvxMWfBcI1PZBqwIZtHVrnHEYbcoXZV73vCXvlQbb3Wx/eQcip/p0v
yFkCpBPxkFiDSY+8haUzCusy8wt9zOOTCLSOLa6L5YBv3Q3a0J4ZmuZByo8pq9LA
Ubkvz1B4jIkKnnsmDHoC6jZjpwtv7l2jEvwpFfXDLO+4d3ptuaQKpqfqnOgtjXzf
zJLfSCuNoknUU9/mBBTRp84WDEbycq6bAi4TXpCr5Tj3S2d7lufNePgFKwBJ3/SZ
XMhaUivAdMus1gFaqjt2fmZiaQOS0bDC/ifuPfe1T7mtenuLSzXoBfTygCeyEK1u
iGMPsvvrkaLKl4gzPzbcAq0G/oCyKQFJkBKrhe8+4EbLYgOQTkpYL6mE++J5nqYT
No6G3DSv0gSuZHJCHwFHB+wxr71Ve3iceS/M8hqwHbndoCykPqlIE1lvU/lPAswh
HMJS8V57Sk5BP2iql0NEahMIhThPlZn2t42LHageX76VVRTaKXah9mEd/BauMjBT
N208u1foIOVZRV7QSGo6n7G9qhznQQmvxTa58pOObG4JBwps630dYqvFHTx19luM
I91s2gSPGJgXoBlP305+ZUVFuSrv7D+LA5RSW0rjfGuvVLVqxHAvtg6WI2OswEST
8OdnVRptdXwNgJLtyLX37ZN6FYZ6qGQy43p144xbUG7e+RVmV0F5R2Evrdg6P5PY
yg90npKl2p82oil5QMlkooCllLdJjDiIDW314PrGOg1UxtvK1M8+ZMXO9I+Klkc4
W+1f3dYQiBB6nFb15VJUH//cd7V1rHi9VlHs0tJls7IRTdOf0lE8SboQ32yj9wFQ
tP2WIpbmKjUkUjjm405ScK1vjbOrcN5a81IAEmO6J3D9tJR+xgEzopcCchBB9xBl
ttNgcC4QBP5T8HBYic4I+GvCKTo/iLivIjny72Yw2u5FSL5H9XEa9mxwZciqiS4c
0FrMsOpzRqdhPjWTQmqJ4wsc3FRarpk432xcs6wF6ZRyPNUTFJe2/MpfNrouvZWt
UezZq1L79Cnb4JuML5EPhqm28p+7rMKl4LdYsVOBG1C6IMo42ejp8N0Cz5kBxRPW
jfyXI59vz/Ps0XM0Nn30K+TgI1rPbh8x2KXlo52SBmdjs8ZX/sinX0WFtKPPZiQz
kxYn0BF3Or7qGvd6wNA3jqOF9W/MW9TQQCWvk6G+LSE1T/sAH0TLcgC7WgYGGIA+
Kww2ikG+s9oBIL9zC4dEN4Hp1qrIgbE/Opk0tp8SHZ74fbb3ulky0pP6U1QYj18Q
PQmUA8kS5sHnK9bTD3dQHAJTyN3kuKtDpEW+SWRT3MeJTSREiyaM4rMwNOvXSM0B
CBUL3nn+4O+8Fg+8r3z19iX6HEEDg+3YlekCpkVZE0EOXMkKKVPcvxdV0AbAJUej
u9iOQemZSiENG+jlDp6oOz3oFf6U+prBvmSZIfEDvcsK6bLcLsJ4KqMB8AbaIEv0
1EifGx+50sOFPR00jTcNYuxRcjP8rhCLmLIP1OWv/i4qbGkQq1CfhxYyPKk14aoQ
jPUy+GGypcMCAxouTQsKmBnR5WkFZese+7aJFFjqIBo5JYQfIvK6zCICQNDHNk0X
8EUnmgsN1umExN4rNvfTlTPfHidFBuFa7NERc9yWExmw7aVQiTt85nocC0DY9DP5
ciz4iNK2BrE8ysf+0iL/5ptYNeARZbNFoS5jt4Pn+xJMm/58yh+L/w6WZZsIiC+U
mDUopkC7N+fJmO9qT6WtAMcJT+l027gwmYmQQ2vNaNXXl+zOnLoxQfdaMOX6Xbsv
ZonREGIGaOc1p4acOa/r7Zj3fi80IQhEeBmPEIiMdbTVig8f2P2Br5V9/ktdaI7J
cjA8R13kNalekhCnyplo6sKmddsCjZA7wdewSkCGs9BjJl3SObaYpl1fnMhtpRK+
qt94h/VskIl4iS8EuwiygtWrYjT+4PiDQsV7ogdejfI3uxUD5UO+cQF/WTiVNXJd
ljIxJ9nDChz7mCmj0nKmrQTjWPzBpRKRkrGQujjyslJaEdnaPBcpT8NNuy8XPlpp
HoqVVmSt+Gdcr183RH2eJIKTXdhDBuoJw32Y5BdqMQn6/mqb6T27fdXEAZ2QTKlx
k6zl03Y1ce4cnBA8/7NdU3mcajJjMyGNpGNav99v12QfOH7mCHL6dl20WgsukOVj
IJuPudNQuNr6XcfFJYmucqpL04f/uLvhnLH+lxLJ6k6HJVV1VXFmNS1Bka7jtZcV
aILNnnaKuAcmz15zB4AmEWzeE2eMkoDNihOaWpRU093w+8nKCUxNaNWWJ27jIA98
qINIqs9NJXXEZYQjOb+KcOIvqsNl2PeC6lKj4zjmm17CKHX0KD8OgqE7qfwDAvJn
MC3Yi1yBtwybpx0g3ZVfuizEZErrqhhD1ldKeBwIRM6P2O7Nhwcv5UF7yyQKYu/Z
v8fGUnRJ7aiKBpLXf80rxgLdOpvJAVazNhRrlRd0bCM8XPeGnilM3D4tnEVaIMRd
AJlbA1dX+DN0f2rbM6+qQ+s2K92aFAhDKxQ1B22PZAmfLbbaXldsS5bzDbvmi4Eu
GqbuBa1QJCxteGXLm2G0O7muUp674iDHg3yeVq20eLq4iquR5moeiAWThy5rOUHx
bWGP460JOk8iXvj5bl9ciLbmvETNo7R3rcUXG5JNt+ImJpJAmCNIwkUifaZQXWY3
2e2WU5l3XeZUXXCBR2VfmwRgttI8v7HUcmOuKsUyEEwRbbL6H7UTVbnRczgPoJgG
XOZD8J3mzCMrEMyZo2yQX4US1W/JaF3elTTNTmHjmcAIiM+05QTFYkbNwVGK23Nd
oMzyzdBGtrCz1TeEQ6/o/HQgPql7ObXqb1I6G1178Qcgx6Nzz4Pgko4U95wAAQgu
e7RE276WqB6I7snsPoel6gOyIHElVX5KBC/2IkBrdmpSQqbuKo9zLhunNlmVdEuH
AoACl8XOj2JKuUvyLi+WX9R/IkIKOpGFt0NNqd2K7rTKYDWJrE6Vxmz57tEt6ThQ
UpOV3Q96OND9x2lhhOx6QFJkPpE/nO6UeBUcmsclOM7nJjbe4amVNjFGlCsDWhhe
UJvJc/gjO/Gaee4EvMwErAT74kDjmjjfVR8Iuq4AGszZiWCwC8yAVQXpNEBo9Sde
+gf9QXFd1SbyJJjTj1Y/yFaKOu4YlLcOWnDtYp0zEXn8h75yytEYWN7ljJc4eeB8
GNouGzQ2xtrXEG7T3QVUDluSpcTtLZ0GO2hqeei3FnCxTD/FaVHbmBur63Yjt9Sw
RdOh8msja8yeLfEXx8XcqwonJ5w0R+9hh1ZrpFOw+vlDJPUZcsFXs3fu9gMBO7NX
el8T1G/BB2IJJHlbFdZnY3R6om6+q8wgUZgdadN55gaSB+bzI4JrA1ZVEHvEWUIA
OqCLA6DAxQV4W4gtho5XA7Zo/TRvUHMBFrIeZbgvOLmhHYglWmOKssjsjHDBSaEy
BqeJwAGemitX2ICrHgfX2uw6NWTl3pXTJix65tiwdVVk0SuDAyag/w60qrxMKnka
QfypSPdDBwpH7q+NkVRpEVaKZwqpOxWfmSZj8IaLI8OomEqYzcwVtVYlDBRbRriS
rmjeGn5xOM/TFSXxtS3yHGhUhIo11WhrYjnNqoz/ik/saBp2D3pngkK453siGSo0
Bpf3CE204C5MrOMh2/tzcH0/cM2ZTw2vkC6Aa9JojsE47slcDCLhepV90nxJuJK+
hqFU4rFjZUAe7Gij9uirWOK7G5efgigOpFcCOwDBGIngCkwPBUF+KdpjUs3ZEXXI
0gGJgQAC+pKM10bwAC73rawRmiebGU431hNRzvX8f1mV/P/QUJ5hjTjBO4iXDmCR
cN4xOh1qI9oCCHvSEjZ8QUxfKVCI5rP9tZGiFly3aP1GwlEDfC78bFLNKlDh33Wr
ZZAdK5DNCxsoBibK5xYGOLZQNWHE1bK0SlpO1zgBq7R0jItJk+BOhPaiGZoMxdCC
wBHa+25pyE83aVdJSGJmXjzKQ71aKrZxath2+Tgia3kaX28iqFbOwPEx+mCu7FE5
RPcWJAi0hJpeUMn/urWepVuBnemJ71MRZgGFvRMTtucXtk3lfYEa12L+FuosRgs1
qbN9rKk83XU/HSJMN2MIwkwS0Yt29iPyHrRWWddC7MNSSNHCS+uHHvf2xLaTDZ93
TNLasIjWAwvCDTewPrEnGI71JXSgl8UeVUfWXGZXJPeIXvWFTajUTkNlRxZAUk4B
SZMGpR9zGpLSeCki9NAJzlIQwrJtPtD6EN77DvvW1+c3oiEncnjG4vyV5yJhAnkV
hxRFlKNYiD4Od3fqQUWpaGn5C1KUjtgl/wTI5myjkGPuq+AfBTwptz7ZAKOKput/
FYhY376YJEKsY7bCjSGiAPdm0LxvEjXTSmVU4MenQbvtWUxl6ouL75cXW/74GHf6
a2Vf3kQVh7CowRrFfkTtRBHWnZhjQE/Ktp8GzqGiUbvmW1KTsgIYBpHuHZtQSo3F
bdN2rulUSVpv1DwJ3iE5fBe3x6LBJ1xr3IQaCjgtk9+3BegCXeE0/3asOf/T0q+f
QX17aTXop26tQMbFaNuEv0tqnLquBQCXOoXW04K7EyH0YolI07kZOocfyEVYZ++T
vJ50wx0294p3Iw0zsNJ0dz0gC/dznYAJfDkjxImy/lPqsYG3AjqAuYn4c/G9Abqs
dzaIzAO3RoBbREsa3xQkTsMUW/ylZT01bDRh6HJCvBCZMcrSQCS7DYVs9DAjekcM
UV+szq0uLRpRS4SX2eLPp8/PO7cGdYqlm8Oa5U3GPrHjxx00d1YQFygHwGbxkhK4
i7s5Dh7LJqGm2LyoIve821JdPwhbYPavFe1IJ01+F2d/qlt9hG9i8V9zVlRlEqKA
lLULItRZKkMLnkZ8IU711GJhdNK+4sgXO/ShpV2BmjPrLZQ4AedlPpXk8nGMld9e
wWPThf8TUcpUS8zXkE31qxtfOFfAyrwH6tyc2FXG//zgbHAmkLc1V8UMOVj8/JoG
Cb4JF9p+3SWHKSzV3eVyGYIB1HGfZXuc94YKphSn3tRwAcSoZTh8kdamBKqOdZii
Z2R1xoAvd52dAqBsAf6z6NoiXUl4VqRxNEnvETqp6z/3ORWGhqyob6Mx65l94eTW
ZZ4vd9UAT6xANqADDuiLdo+DR53zyxMhnlx3xX7gzVDRs5aoffvbgIiPuHWRcKvi
rpebGw6IFQ0uI76Ukbsf2jWoCVV9Rm6Xe4HhBITyVIWi6jF05Ow+FdMOxk97Wkz1
nbo9bM6NZSB4NIvRieEur553+l1WglN3AIq3bcu+7HBJZHyB7RYBk2zjnMWO4UZ3
Ejj06X0mC+9aOVqEwihnk6Y83umMPh6RX3qrjz0t0drMLYptU1N1l3mqkYOkpk1j
Du5qtR7PHkkczFWktX8K2x5oR6V6NAOusIBs/kEwimUfOglWAHkvwEMuuvKocbLp
epXoQt0m7TLoNRwtgroRnF/qK066IMuAKUA1ncpw6LJ7EQBNPfESXdDfnly7HPyl
TG+FeZUNeB2Vy5eu1E1MTPRTeHDcEbt2GoFwo1CgoboLUF0qWiYGozd8j/l8YZ40
l1eCBvakpvyXhTuP0kvnT7G6V2vF9X4feLEtzgdSM9EJkqV1zL0keWK7CCfVsPXW
ampXqNApBCutKh78jiS43DB5C890tUs9qUbWwFRuX1BYoK++dlOMMIxQQD6gFm3X
cRSlyJKrfn2gvc7MGddcVJxxox5mMH8LOYp0MWmTK5gBF7TSit+6axGc8gvfIfVR
Itlf8WwjzVxQ7k/Kl4+oAJjIhQcomb5OQgsDIwnOwfjHxy65CppvD/9tyLKXW0sb
7sJSpelwbVklTa/8+8FspFnuiVwVla4ORcaYgcyCHjfo4tCRG85+JEvdHQ200yET
JnC5c8uOMk2L0n7ClVM9kL7YoHTRjq9n0lkDiAr5aTprbHDWllNGny2kxfKe1vAn
nqsWizorb7HhO5MWvGe625m/sBg0F/fAAQSdu96d9OxgtI5vnMQpU2KmfT6VAhhL
UQ7kDIGy+3akgDVmSy8hGhU/vOKkzgvjqfSuT1vd+rBiuFOGqdTOlil2yj4D9z8K
9yWCosRLsqmK/JsQkCgHt78/Gzjtei3pAFNHRCumZN7bVgThhf5FPOu9HkI9VH/7
5IlQvMfYwMH46q5meO5qFO/3kGyoHjWU+skewZ64NspoaCViRtK3l9BDZ96ThXUA
xae1eYVKZhYImvxpsIiQJNXF/3PYgIBHTLTzRrM02HanhZY8qtZPbtU32k46dWJF
wT1C7+IXqYBPQdPP7MHok9iReFC6L8sPL7SzjMnfE2TzbRHUtgDFEPyhuSMV7+gn
Xrrt4YHuJAqbtE01Vg0zZ/yoINg8YOBirMZfNypyke7zk9gwLti+Ix0R4OM9hrF4
l7q8SuzVp7BpqG6KSy0UysnoBhtwtP1dF38s8e5ms2kM6TQTC9JqsA+JgRMngtZK
XV0Wb5TYCrmLJihuYlTvOBfB0pSDB9uMf4SUpxOOVXCuujGrDoH/FnZYpW471vGa
ux4LOq7ijAVQ4iIWByz1WH/Vfd+Wwujr0KfLsZMGBacL0rHPe0YNdr7sW2I+gRf8
lP0hU34s6dzllGxZZMw85EFQKffOzqr79+ICeILwVopTn7QEfi1QZ0jfWFJbr0ch
AHruMlILhqpRt/FAtVp8Ydck4zaJl7ceL1KO8gy0Nmw+lky4m0Ff68xQIePD5WUb
GaTuHUFj4oe+d9fBfLGn3JfW0EzbktXdEa+mjqqHVDAX3rdX84O3YAeX2J5PHA8s
MTNrLK0XqdbpHtSo2VRMrF5/gCVbDY9nt0AlE6dQW9BaI0/bPqTWlnTKd8TLTeMp
PKGjxAnlzdHe1MrkGChwcqFK2WWw7wM16LAhasI8uhQbtmTirT+TEULbPwyCFwsw
9dijffo07c1P+DOxw3I83tYTJtrzml+r9dRiXk6j8GCbfFq378Xep26BOPQuR2sA
2/Gux2fHugB5eYfkanFhk0r8hgqIiXaLtUWpZWBA2hhJ/1DS60iZYL8deHkFHksQ
ZGD7C02ZKLNR6n/uiPBvnOwzutnKcOoyu23zBwDDzBef/AxUUNmojgKzQmmsYzTX
1384G0AtGWm3L8sORvcMcdy6HIa1AkrO9fEbuKAmz077LvMX5rNZbdiC5WlKR+lo
9tAFoVUTF1BGi5ikrG43h6n+XFEJgGiCXpcRZYgYqGe+/mswR5bFHt7Q7SgRDfKJ
1KDPy1I+Ma8mjSsYANGAjtOtLP1h+rzvcpnrYx3AvGwVGf67jq0yvb8tpMlsgWsJ
7/r4DmEWk7IomgIRj2R+UoFc2U/qy41L0pwYWi5WmBWppavJvPduKisXlBuGwYAe
H22zXDsoCxNvqVzObGmUuNjrSlTefsG8zzDhCcvsnpnXoUEcfNapGgQaUw63UZHo
J3+5QSp5pB9nqStK+5SAC8rVjTjYxTdjexKc5Qyt65u/5xYGZzheiQiEjsvKPXlw
SObqNSffrri2fNqGl1nFVn7fH0S59dTrRPPeMDHpoGc6TCwgKggo/BBIktwAHFcN
brSIcVuU9qTMKTO/XXbJ6z5p85gMdDXreHhMvNHtk0ztcSrLCzzXJGG43w8Zv6oZ
ffKZGLXBaL5pmoMSlbkVLtDzosFeBeSmayeckTb3fXKPTuQvQQj6q51koNftXGKR
UIgjQF/uxtjBCNqMZswhpbVIU6V5zcx0YI+1UPQm1cW1Uuwm1MCWjXX9GWV2ZK50
SFUcH91zSJSsrqluLRo9fH8U2PXbZsGCvfWK/MYp3Y5Vd+K0T9hGueFupYvz51BY
kHTRB/P4JaLRBVcXXEiux0LWtXJwbuomjrjnXFJePwDiea1fp5ngrHBtszo6jitz
zjnW7MnHyqBUG/1QX6iHd4A2a+Fh2KOrap2eKdWow6fiScWjbGQAwgmHnndimi7H
T0IdBmj0xlBQBt0bWhdNZS4thgj9KbQ7FzKflx3Y6ZT1eifsvUacszeFeuWBkods
YeVSabw/9nhScTxgqpiIlOGJtqHD6QRcN4Swus7Dsw7H08fbc0ug+84U+xLz4FaB
rGvMj5BpkLlwJTSkqxq4BBKiqUd0dRdihsJiZyqmv2ayntm1Z/x73QA4sJFpGgSG
k+APCkZ9+JwpPJ4AFG7CXNxxNksHofzb8aJaL9FkmKGQkItbAK2t2jpK3hNIgw/0
7TMGDDNVRmYMId0AQW0yaDsMMWNpEXYupomG2y+HT0sMWaFn1gaqhfO18hlKJLHU
fvSaWdqK1O8izEBmGXBKSC7T8Qyl1Bc03TXU8bY0KT0/NPVYZsQSB0v2+i2jRuTK
c0GwFF/QrYUD9yz78LdFZ1y6C85XGzfLDxr5alDhXiw/kzovehTxwU6xFoBJ/7BE
rmzduFqw53CDEoaM/Ba2qRGev0+gI1AvCZELrDxTtlkv7ubhNYtJV+sQFbjrqthj
bc4ybonLT4o/enp8Flxld9NoAU2edtjw+wLUUVcpbJq8zfYg9s2N6eYM2K98/KJX
Ja8JdZnZbJ5lYjDeRqFMBOA4f5MeGI2GywR8Dpmt5Bc55Mykw7fP3cbSlDxNe31m
GaTywqMWNPdKY6PmFU0Htn7vff8qIfWQvy4kI/BRh7qFN/eYqPRcxj8QMeHw8r2d
88Ru9DGVHW4z/x0QY/sKIf7OwzjFP4Ayyze9vazGVghJ74dOkRqccGzXG3GT0lYM
VIMfuhtZa9ndDPEogBneWBi0gMKfZ15e8sgisxpm621MdJ8a/5O8YVPzMZyRnX0p
/Hd4f9DnaRMuPABqKpqvnuv4kx3c4eMQWgpHR3pO1m6TostExjN5GpnV0GLFybS4
S56KLDsPjd3BdcBru7zEdugvj4mMPolBr/RnPi9jdUdYCWU/7WklsI64ek9BjJE0
vFFi9WY1FbQEOVGe/cGB3ZNTeaznw5h6THc2EoWKjbHu8vlX1+55H5gPiFGFqEtQ
kICfSipndZrECZHzCFKWHQwG55nYWlsBOyGfX7nE86mhwtaJ81emSqFH0uH/pU7o
WbPBSWWcsR3YGTXaLSTbVDphCNAtRfhBPok/6KZ/cayPfH71XoaCiLE3xdPNho8Q
EACnL+xEFrp6EzcL8YT8MPkr5dINA3rX03+CLurBvBJ12uxXg9qrue7VXDoXbGdd
mp0L7WkP2tf2G/60hvffuzsemQpJ85BTAk/JUMx5Oppr24NKeqXLtI5XFF/UGdaf
kF3slH3BkeDwuJe/GG5/2NMB4fmxQXbWlWLc+kT+bedmRNYhStYlgMyuhyjJiitj
E6FDgGyyDetZv/EKD9acaFIYa1YDdvk3ywzg6OY72Gtdv8IVg1BaQVCMWkwOhVfV
OCM77hAPAjGxMYTbNOue3N5EJRdOIZS/Us7tizXOrb7JxqiZFKRbwMcLU9nIOEzb
faznZuHX/8bKopFM8XeTQ79svqSi7uOFv/GnpvImCcxiwc8pAkF4I0pOtcbFTXhq
Ean1vC3nBWVrxvQKdkULad4LMyNY42ObIBpAurdXkNQy9v2W1oIIgnPFOUr8aIrn
hv7xGe8uSg+PfYKMRn2jPQfqd+uiYMq/mSr99S3heyMynhgUZThWsLm4k1Etv3/W
oge2/OQhlZTpiv+O7dZqEjqvskTeZ+ovJBz8Ynz6UDkCLEQp0RWCsjNyuAnOSYKT
ducFECdnH2gN6q5VB+lm6XW09151+3mHczPW/5cCT3GpjbLKARtkoDWkf5rN6ZgK
UfJCfV2Ii3w4ggKY9JvazDsmwT5a9gXkb9cWAG81NNmW5iqyv6Cq0vC8IZ42v85D
3Q8PUnU8jawzSv201m6GckKt+ZzUncwtWxJgemJcc4tzYhZt8oImCWw3V/9z+gvs
ZSlcOeUzsdsTljrM7sIujClSKxPD0dz9ljNrn+pG1vh3mvXov4PTK1MuvseFHcKW
PUszh2j4h5At8b/nE5GCGfm1mBqPppmM6+RXX1ceEqgdps3bqRZq2q+3tsAzP2HG
gUWhe1Bd8c7Osjj0KaG3L4qN5qBsSpbifyZVTED9OjTgbuKDNtFOY3pR2+gcO6gW
1uP2rurPkgQ7MUxbo1cBwHJ3ADaAOhd2+2ubnZgO7N9fPxOU8r4hjITBR7H7+0Nz
1Srdob0cW0ewJIltnxfnovW/UqWCDSbijWwITcDTdOgDIYY2Nnk62TIS1JpG7GMH
yfuZs8Vv0expdbzaUuhmHc3USF2GrOriij7J19900Otw1T7bfXtcWDYjmKvWlIYR
a5K5genPhTbo29afUkg/O2jhhRLioW0JhsNoo6CH6XIKL2C8Cr7hhx92HRYGoGZU
GoV2MiOS7epX7mGmr17YkxXFbpcue8JbgKRtUMmTovy5nBG3WOtuC4ZkEtHiENkm
w6w6o56eTyeLxewzzO8V0gIX1azJbh+RzJVBBYcebWyiW93bxe/JMphKtvb2aM/S
lEmusyj0KIxUnmxpbYUAl0noBLZ3wAfxt+U6cCwLw2nxPjTx6Jpr3H8r6fRxd4QS
rYj3JwBxRtBtYhmFITEYd2dpImSGYGtnTjJnJg1CwuA/tguxbficlKplrRnVe48E
JOHqbTlAhL96POuwEwU9ngfidDUG+GkyhY2B6ybTXIF+lNKxj9RMup0F6SErM4NA
KfcjnOXRwoyxJJ6qJ4GbGJ4uelVcVv17XPqP4IReJQVEp56J5rQGav5RhvAxkN9z
TlbyoaSu66d/+Jza6NFc0vte3bpuNYaa6kq5HgUCkKOZpvD/k9fTTi9So5lk5PoP
2RwFpbp1se3To8QIEQzfWWdBNCexVDgSGzinUdRB/aHZx03I3AKwgI/gKmwWd53L
qTQJmh5H6ULc+Ou8dW/FW3M7uO0aR/xIuliFZJdNkQKRuidP6ZUzHqDIqEH6uv9l
JqUVdBMO7eb0csDC4grfWO+Ns71gkqtbeT3AfyZIAf97JLkyDq4axJsmyvC+J1A7
WZ/4DxyBt/EL89jqrbzzuyjmzoRYmmV5CIxlDzTzOUuA2VoAEt5y5pzvqbo7rhbv
9rdglBTRMK3u3e66WmQi3SexWtlBbbPz2giM5/0GN4s8GDSHZEhqfRK+rrGjrDre
wAO1Jqpp+nelw/fLzWUcDorDaiAQGQj0EGv5t84AcP2uRvP7LhxlILYJ4ce0aRDU
6YRprTZaNyL4VjqhMsj4of5vr1MyFxuR5oIE0p+ZVKzDae7sXgSuzE3RoU8HcHy8
fAOM//xJrazAtNY/sRi8W7x6UvDBDc35qb1MYd2dS9saUM62dN0gtuvNyxbDvf0Z
Cm4luxI5NejCMjswA9uJDth58sNbRm9tCyww3C1LlCHdvQ0ht47zPqOUu+KBvBCJ
soFJQTkjsBvlASIX5bLhmsGXcS6KEE8LGUMQGM1nO2WVAhOhscZ6T7G8gxNCmHTK
fEvGCI2vw68EH2TOHv7tKjp7kRhz3n2iSopz4O/+8+fgxzGC3CygDzxHIFcnotCZ
iZnmx7yqh4KuSxlQqcX+Vnx56uyY+o5uK/xhgLnNugLDpBSAh8Ei2mDwsUaXD/pz
3XPE4cNHRQrpX9PooO31I19T8DyWvyJWE1imEEQyarXB46msZu3hoOyS1psvpa0t
jPx8q77PzhWw1N5ka/WLMJooOTIsCEpGMP0LCt1CZPPTNirXvX9uFE4A+yn74408
HZ/oVm8TbDKGnv3Ovii99NYLw9iv48JRkh/qiwf2OMHIl+U+YJorLjECkYznQtQ1
OdCgHgOS+FFB29XVxQ8XfQ3lTteRZUvqG89q/NOwMYqTqjlHYVV5nGVQcjkT90Yx
7CLTacm9u3i5Qlx1aZTF8vfS4A5p28TVU0w40Gv2jIBoOBxesXHDFjD5A7V/FV/i
nI/g3TXALUYIvxDxdsycFUUTrl2wUfFz6Yu+zS2HKTzXQ8oBz2Do+M4ejViAonUn
4N8V8OrH9v3vmQIdPl0pzFvgNZ/3DMz8kiNizF+/ldG1Bt2aRGW0sqMMOLtLwBST
+uL3XsH+ly4XMugaBRfarg98eXnhvpVzEB17z6aXHeREcYMPimh/HNxf4VZbyUqz
gXxrSffxK4XQYmVKUAUkTXOxIW1pRUz3zZqfzv5wXrNd7TZpOKszfBLud8AFXcfq
BAiJYxQPc/vjUcs/a4D8t0EnkGqToxFD8KXA5QzJCT1D2x3KwnA6aCqKdG698ssu
o/mXVHEu8IFdylJiy9DatRNs6HHDU+kM5gV6NqqdGpKrn54UiWlqFb3C8fHt0FDV
FogmrbhX0QpO7ddKRjjUKzljKOAmhlYh4VTGUCEyv6kdJ+IyiHrAzSK0rlrSJBDG
2XbzGQM+Gmc/dnYJRTPPv2H6BZq83WJLxMCZeN0YIfktMX/UNtlunxkf+ppv+Shn
E6WZEWGmjP5dATOMIKrkUlXrgwcP9bEqaFc+pDui/+qAl02iyoa2++XPC3oka7uL
+obk7xZhmorkuc/LuHLPfDQOBDOiVcHVvjOn8L5m//jiDMcZuo1h66zxuJu/4sqd
KEUv+7I0pWqpI3gzKi2YnIi1PvRPIuFLx4D9hyY2RrZ3HnKEBlN8mKGEHaefZjBi
BvSK5ZzWQow4Vpd2Wf2J31WMGauGcntF7xPk/w2xWky8ryhpD1KtrZcK0M53tQmc
0Qmi7gv/l6h4pgM1+y+9ZgrdBqlYf8mcVNqCC6ij+D++AvtysAVDsaGBKqByVsK2
QcDss0XiOnS89k64KGzjyHIZ1uzdEC8gn7EcsDuGF1T21UQ4UZijh22ChYTqBtmo
3BTcRRkJ+A5U7QMAQ11W9Y3JaPNjfwuMLdCUNsN11ldBmZLxR0ZbgKbzEgDlcbZF
re0uEN7Wma5ZfT5zJqs8zRzG7Lfsg6yO9vUJdmjO6wnsOYk/alPk9FwKhF8xYKiH
i4wa9VvC7ZcFgnlwVNQnvdNLi7g+8bgbeMzkj59P8S7HUopxw2au5WrB9GajqXYm
JxD/NpZs9TFr4CTFmNx4rQ56qZIJdfAOmJig9TOWJiYiNOfVXynVWg8o79BIiaYV
N9uifyQwwjio6vyKP6ohr3kZdw9FPvmyFHBuWgDqQAkiFqUF3//fNUWS9MICOoM6
myHcNhKo768vfDo/e58mC8YhcnyTxaOJTsn6SzQuulcXcMG9nMJXfqeMW7U+bKLn
7TMVHM/KFiM7KFicr2htTAxA8NxB5w8JnRKgYbnwJNFPNQl1syOBOtN0qh56Cac0
0e7h2LfJqsCF5yzHg2dgu30I7yvQPpuL7cajU7/EaGWcRWYGS+oYUabfnkVVImb9
H1Ys4psq2nRh6B5xP/H4aUfblnjueZ7IrT4eo2sICq2xuUDtdlTbWMogdYy+0um/
lPHfYUC372IgmiuDM+Wu5GEfaeIu+PAXmJYekg2/iir1B0YfWdFvP9yFVSksC13H
WOEQhvW9JDcKzSwnSyhrGzpZg2Bz+IcL16nyCEV2rtakz5urRNwybuEpRZc6IwJp
YD++2GSuz7IeTVjcBfwwGaY6RxPErLjmV7vXgvynJjgt6hVYsTcdySrxkTEF8l2Q
K4rNhZOjL6xIWkMLIuYOh92cqNKT2BszcSJ8qYxVMJOvPplFFV+rlfErAb4ljmYx
ZQV2JPcmUHKmEOFvdQMmanFgSvYcUYEL7jbnY4bdm0aBdRSMngQ9swVMxDlWhcab
7oBulduK9iXSudRdS5oKKFKXJ9VWxewDagskeog6TYWfqZzznQ0QFnXIut4CBdMF
8q8/EL9EXFWuDPe0oq7ALeol+phSJY4DaT2xJojOdwCM26eTVPuzK9j55zQghk/U
GiGca3AYHiPWICDqK8R4NUht862ji2mgqmyqTFRJK73YLUOeCJ7qM6JnO9HB2AVm
7sJBQQdarIeen2nrwKmPzvgIrlmegdHeyRL4rKxf0pYQu37s7K5P+DAmqA3tPt7S
KvdP2XJ7kseFyJO+GzsGgiKkjL06cuzTCeiIGVfnirmIR+7qhu+VpWk6f4XmDHkE
KZt2r4GoODL2y12rQ2Y83SUtJR8wY0saVCeH6PGxkDXJsaXumoSWVuXgGbGhPIYw
8wI0BH1M0RaVfttBhSBh2EwMslkhES/xCUTZHOXHL/CLKYmT5EJqCHCqkvZC/ori
dba4b7yaa3XgHe3cP+lkiUK/DByUrQl1mt9Fc+2F7RJVy9ivQVr+pKfXrMlI8q6U
3fX2OwRMFPLgbcmtnuZYUMRjAAezAec3ONtNrSEl3WZJ0R+v9nRrQOHEpKQtc4Aw
JbvIm4lVKw4RkNLtzK8dZ9vWeYHPE0IDSjmZrLuCH2SWipcbt0W1QSIBJBo89NQ2
rkoCWUWhZQoDLMlZCu/7Cl34kZH25tLeN630H4MgtBe6EY2ir9Opndf4q6m0Rmyu
i+5st6ivomaBmeg0vC5evnfJ7bT9xGVoAHXS6zbuX1HMrzBPjjxLdK9RZ0nfvzQr
lC3JOytZDJ42K0cDhiHjmYcJdYGUXOMycQM5SZVtHts0Nz5EGjTrPCCyB4wRxuKk
RVkwJhhURoqncb01qhGpc/CQcqYdoTWu5I+RS0abFUBv2H4ZuQCSezMIR8ehtPtN
QHWbgt6XmCUnY7ZMlwgr4ljfI2d1x87lRJQgnPJea5J22oyaqD6k734RB6x9kYgv
EnYg//OaAyZaRdNIlFquZbmUBBvEbU8twBpDIfJpdt/W7AQwZaT/KJ/unyjaPHBM
g386clT6AetThX9bNP7M7tMOq4EJJvdPMplfQGM8Nl3y+CpZHRwaAjl+jyDsDyK6
1bpskIeSyrgEBbHzarkXnO4R/oDH4//U4KqxQwUJ3GKWeMxwORR69Ekro9Z322Hu
b9grE3ZCZWCOYf3t9NpoBhTyJ/YwloQKGzjObYEn/yrFvxjauFO55KJuw+s3Te3X
Y3Hq8Xg0fjdw2n3SH6sxUNFJa09R1YfOGmfNJYD79K2xkxpNLsV9CvFCdGKwSDQd
LaetoOJUVQFoX1AYi4FhuyomXNYj2LO36v1AiZCo+4OzhhmLBu77smeUGV+SMCj9
5n+9mRqJp0gohi6BAUJIJ/ueie8AymsHqqAgJjv4AbzKA7tM/FAOwXILPL1y1GvU
sGvA4spgT0bQ1F7blWxnsTZ+JUKrOTQ7TAwae2Q7pygAeI4xzUAjC7jgf1Z9O8Yg
jkVVFr0olD4fY+czI+OYd5HzkRlfkaD1P4l3WFl5Ex4PJEgTRnO28j8N4CpzJ3a1
sZrNbbMdTzKLWIw6/H8egLpotQp51v2gDswoRe+KcPvhw3P6QGxJs+7OpFUTvJ6b
rMQ9UKfRwOgo3iyFBpKXjZrxoZa9R9LVfE/N48iJfqIR64sZU3hj0v/r7tIF8Zmt
DVcedkBVpJMjThCBxwuEUYigOQxBzuTp++5sGJYYMFQLuZfjsoHYNmQ7GcIr+nrP
92+Kkkv+O6hSuafW+Vt+7CkY5iKs/Fc0pIK2Gk0wZZITiTX20F0bEWKiBI0fekEV
uLNkYJX9MqiVP5d2/xBkNWd18T2VsrJx8n9VGo8wF+6pj9570djLVLjVFuGsK6VU
fs29HXa6SaVJ8hbKaYYfWDVI0E4UkQN7h59pZGJJmiUf34CVn0r32gIA+nnnJg0m
y8A4efq19aBCmf6oTwezQzSIRxWLyp6pFvW1Xx/uMkUZ4cJZnbm7iFvzlvSWNRw/
yZpHMg89IU1CR+nxd/JkCa0Kv35JBCMDxNPDMZUfViLLb3eRn11k5kZJ78qeE48x
wmfB0j3iEsZ+QcN+dC1e8jslePmqQbrQ4dLE171d9tXtVObXpVJiQD5vsEtiqEqC
VKOdEQUfH+plnZZi8vRP+bZqf71xwe6krXH2D+B9CGyLkGDdpqWITy8EhhMf3Jxb
djYkK3Q+k1bmWCOEychIS+ApUGEgYlzsRNOV9VKUY/+sZc22rnIDVYeIMQob7hge
x+j/YdTIFkccEJ4RdqE2xsZ/gGj4YpqQhobViUCzdrFyL+thDKowQv8QTHr3xXIz
VoJlnVzmKBM9BNN9rI7fb7ZpLOuYhXHJ+WlBtiQBYqi7/gADmN9/jJWFMz/p89IF
6C9+XBatlGafKxPf5mKZ48nH51CHzFjaxua4lPF24svKDM23Uobt8aOsBuHulkhr
qX0k5kCyK/SIRu+Sd/NerlAO0pspMMSq5qBFncdpNyWGkxjhiwm4W8Do9T0rZIG+
jsNGlwjUK834zOzcBDbPsIPhIXsurTDfgPwo0ctXhnj/SrKb4jty4AdFvxT1jeGb
OCZS6sfGp93HhWfV3pH0WoX6YhBxV86+djKkFurIe2fp2+CWfHHlJ2jAAb1Z80X3
nymHjk5P705S8/Xeakry+pMpYvATah8m6s6vxX4UhJQ0vQjNgsn/hjMdOm7eNqWJ
L1nSdPem5QNt1t7QfFzpnjMliPFKmy1G3I8mg22q/bbvix8fRJHOsTVrNALugfdA
iaZXt4OeNyfIihzYqsXlD2I4l8Z23vPRg2z/taXOu4KLA+/rqX8hgmrQ4E0b3KYq
v4ja6cVSPY4ZMpZY/67mxNYF27X3UvKsbOyYd4CEmsGxvCx3t+xBwWo7V0W57201
+wotD5eBZS0Yn9o7+2tunzwiVCp4wX/XN+/KbbsLsJQmFi4d9/L3O+L8s5jKIwqm
WY3HamFTqy9Zx8CTjjeRPs4CXeERg/JRw+ToqqLyF8LO/pnv506brhc3Tb7rrP7T
H2m+sGMIEIS0d+IdZh7BAmXwrM7eVGCXZPU/jYZ5dU6ELTMiVeg5b5hBK2Q63hTo
BL4KxdXB7bOAHcj1YgCGwukuo9quXcZhnAiirEdcfJpXroH9rtqTdv9FBfZyJbk3
BKhYpjRqvgaMY3rHQY00hSVNJkueqhtXj9vg4HkYV8IGAqZ9bNv/8wTZT1xi3klt
kL7qY+62xOc5kuXBM2qhs7AUlCDywUoX19abTt11ZapWMNkCqKCfG5nejosPOHfe
ZxUkmFv4fA/CHr7F84Q2M2+h3rsTveqDrXahDW5vdgN3DLWun/dXvS3IGMJ4PTM1
PzJvr90lEoiIT6SpB+t3qJOkC0XRLPH8/SnHVATiT3vPxX3QBdVzwCM6YCRZNH3o
rV3Wm728vkhWcC9v4BNyHSMYLAQMw3qd7o/KqY9/Avv4zm1gRr9K7rI2jGbtCw4u
cR1TP/S51M0ZU0NDS0cKAl0GiIAUCpZgx0bD2gDhtPimN/R0ntYKx04dtnrEXSKP
CfzwowZNL3tqoMpprEFiQHJSMUjr/2VvOA1JwPD+v5iYMUznusij0OxZ/J9/Ng9g
pMtlV1/5EOf5VIeTl33BwZnTiC6KYkZY7in/1tWnZUM1fjT/JRaqnJ8clqzqBBVs
jio0h/PKFfgCoLi0ZENm6OF9sRPBFSXU/a6FqPNA8Z9OYNTAiss27WDcogJY40pP
9GInnNqDgyJwRb+qH9PbTRzQfqQBL09ORdV33gcRw1vuGm238CH3WOTDKXBR7Sj2
Y+5leqvy7iDiAm+xWDOEHytaGZmRWRujPontH8QZ0dmjXGpbzIWxEI1QObWQHRuU
hf/I7CmUaKjy+SisnPfYkm24RweI+8BJk6jxPCM8vPy2IWRLfgLcdVBrEeQZkS1X
b17wHxkF0wDfojpwFW35P9SGW+FcvEqkRQDofzmFwz6st+N0taCrHZDaPqjQc0lc
vBX9nfPigRJFSfIixZJI+UjUnhJiseC9WqWOvxDSG3y43BvsKSYBFtWJnkl0HPdz
/BmJiUMbiakX4/pqSrR28sBnihyz2XBYw37CZMFDzi7/BIrgVxvq7WjY3GsUjZmQ
IOImY+TIgEtHyJBaW9hQobYorBlOoYoKY4yPCokCFAG/EPWa4yUYOW1ZZUDuJq0O
zls3QcxUyfBy+3/sTGPRPBJUuhIBaqW5F3oiuOXk2V/fbYWd/p4pPPbxXEybJ+lE
AdUliuigDW/Yb0t4pUW/3QXgRvoqtBP19IZTyhDBAupAEKv7fm6u+fIIyz1LtHl1
RGXB6nCMcSGUmJB2Rk1+XdPL+R63VfXJh7TC9yXju3Q4uSuSuhdRM3Ywzd81Uwzr
as5UWOOPXYPtR+OTc1szIjCs1PSYYfGcg4Nhpex8VUv4728wyLtbLIZAdcEaw10E
4LWx5YQ9lHRwp2V4Ok61T8iHY6loOUmXXxhNWeI7aQsb/dGutIZbh/bH1wlSpdu1
q3ZyPmMkEzo8e4IQcalYiuKx7yDqIypkyxL2bdw0EEb5zkz244X1DZL+CtmMvn9s
NUFxcDsmi/viWK/L7i80v2Pl/K2fld4GmtQNfHL2FGhsmhjpizy7Jub+Q/1OaH38
maGiZEr5fmq2MTqhoJB/w0wzWZq7HJwhcZZUPjbFO5Hff3CEAcPzhA7IbFPZAzov
XUXxv1m9ppdx8hQyrQDGq/6W4fC9cxeOLmVrDzL/aUUUVTpbekzfW/BbYl1HpBdI
8eipOMUJLjdh26V6NcCI5xm5+ccA6A0K0Qrqc49rD9lN7z2ba7saV9V9e+h9Ogz2
rYREEKiRG7kLGuFcuirU1NCxpuT34XoaaHx5OycOH1O4q6FiMPkup/4sryPnAVKc
NNOw8VtrNWQTyj+mQIfe1NdfqkaWDo6dB+cn73jRIw7yOQYHw77nkG5OIOtPD0x5
qQIfCk61adO8c397Pt6uXONki4rILok49Y/0UZ3n30buaIp48IQ3GVlsvbaAisV6
bqPNe44GbOfd4wbKbT2b4/XeyrgaCXBduNRV58qestk2zga4KIJzgBn1aLGyw6m7
YuHyKT/M0+k3kWitmOTpr1N5wnS+W/N1qoi6/FqukSIKwLLpKuVxIKaL0yOQ8NWA
TGLmh1zEMV1RtDhi15QAlZhG3mS5PbWoM7IlSSnuyp6nzLaNWkwc1NZFnQ/PML/0
H0il9KNDEZNL4OgCQgeXIImyvmFptzTicteaSkJOQxRwjbPY/kRPrxdyDm7uC0md
GcYkkT0Qgq1fMb+QSMZF25uKQcKDssHDT668hM/p8abaYfkWMrReAO+j9vXVjRHc
uCItSDUKB7LqdiN3TU0kNgI65gOGTErhUGlgaEBlQNpVbODo8RhC/Iq6awghb02r
NLm7CNPiX2kkYrpsUQ83W5PG/pQCy5w8JwUYJ0c0jYgxY7TZ1zfsd7wThwNAd4tt
FXrhsvff6X9mPCkXGrRm0wYlxDUpbzycMRTTc9faWwCN36/Rr6Upa202RS0df/Zh
4ob8FmUPqx1GA2ysCYq7JxR3IMN3ExxUldR/zl/ubsmdCd5zA1BxFoukQc3vAvXU
5UehhbFHwX++2mMGHnWSdG70iH1TdtFW8vGGL0DBtuWDDImjW7Ys+ik83vm2Wd1T
ZYW/bjRjWworp3Au/ATvpXwgQ1oxjq9TuDQEKfCs9ofY3cZtETeP1xAE2rEMAKjs
1yJkA1PNrw8iLxK0BHMTlorR/b85KmFoyMC9kq1kPzmOJ2TMCY5LjVEA5leJX9R5
MfXhtxoz+EvsTHLjzmMeBufP864YgFpu4ame5lcTFhq6dgJUFjq+0U4A81GcR+z7
qauoaBep6ztRfsiOyWArQtpXxIrjvA45Bjhk37kmHLhheXUD7UED60oJLRvfoJ/3
oZq6vtxyTCMHSgpwzQRcFxU3JBgnQV0QBF5BgGJycGx2sil6jYJooTxD9YacBKWX
atAeGOxdM2VwfrnryeUXdb9n8KOLoIZTn/8kl3U789fhqDrW91NT1xZ2X7kxnxZ6
kl1LgoNz3tpwQ2jrFNiImCA0R7VjSJq7GAAAPVzemksGwqyxNj55zkjkxda8TaPi
wv821yJ3oEATTnMjYGYvdgCBC+lppte0zYvPz8cF6SPjiTGHe+0UwCD8UIzxVCKp
bfPl2WBVJTqVhOlUqL90tn0B4KVluHTF/JVVteuYJVT6ugXaRUA4aTq0hnUsCd4j
XArz6Z063oU2/9t14EuIqeEuZaHveIj2FHFUNXpG8wIiTnU9vIkwDjwcmwbGY8Tv
K/qqs+L47KSLWOdwAqgNKPmwaXoYHg2glVuFriAzWqqw2Hxiostu11XDNSnHqfEw
WVt7vclMk0VeWQ5FWC1Dsl4XTCTPxi3TsvuXaAXkLJdPuiVeNAJINe37a6VhwYio
hShAipFgCaCcj6kPNsyR5T9ofvwivdMT8SibfRWMf5m2wmUV+9FKJb4VjbmP7n0i
XCCt0tP/aChQPQ/GOak5WOuhdRVGfoTClRWqGNejqMlQ8A7u3LUF7Zr61zPQzvLe
5lk3LaEuyC1HyVn9lrws0OG/cJeLvo6Sj8shWaUKJI8MXzSAKcbYMyep4o/NQ0uJ
6ORCxaFB+SgtQFQaIF0+QAJ3U62XZJAvDzEQKEVeIlYC8eaMGFPkhFdBHH+dv7iw
mFsHi/jJznLjudJbze2kkpQkcR6Poi9blkZRg4savcHYcobqphc6nkS7brHyocsB
ApxAUrX5DPk291FiK07WnqHdvA/ut76tsG2whNcM1QZjcPme+6g4uN5wVoFKEDiE
/2/QzNE4uOxgnnYXhNA6ZWPMoeqzDtrJua0QImTTfgGhvXWq8QSx5XLbt9kbgQNj
EATU7+jeGonEJm533HuCooI1Pvf+PbFADWcvPKprgGiwD+Wb+2zdSWf599t89LoA
wjzKi1pf3vE5mONw9D6Nc9tsh4ChxGz72JNR1aYhBWvKZk/luXJLJLPS7kMwEc0O
/2kLKPDT3zynDTZmxEiiilUwr14ym36N31E1QtYaO7lTPIpul5MwNl0wSNEeFd2k
NIVnw/UST9CPibsAXEogZmPXxiZnyGi87DW6BHQ+RKSXHOmSUKwOTEg8HN8KIFKU
FwPONaTFEqIGlDJ879zrRk1Rk4jVLr/3CBwQsa5dhBhD/dQuRCcMQnDON46v5Vno
i3Yja1q6Nmva1+HpFIDCXj7bHIqT3anVhhDE9w5FZ7E3WV/k3Mm9PUdKl5tMq2hT
JenvpLImrbfk3hcmZpikCxzjJL2OEdaObIjcXUnviRO7GuW9D7gV986QRFa6l/vf
tf7Gow1CUwdyUzfJESvgR0PnTs7WO8S3v327nrYkQUJtRaZFVbSgY9dlNSdPneSe
FWZiao02i007sC5IBY9xwN5SQtKxVXzy4ldJ+u+sv9jE4gtVrqNcqjjoW4esLCLO
rkJtYAfXZcOf6l689fE/uGdPBLE2nlTOCfuuTflS38sWVcw37ap72KOCLle1qrjd
mXve+4jc8lawOp6g3ZWz1iHemhwLigb9ZL/fpnviZ1eo/yTrHEIxJC/Cvi+fuL31
LaJMI/1ORN29kOiFPKjycEioDl/8kmrncqRvIHi1Fn0BUmsl5aHiMGgUJMzRVQL1
37MG2fdDgCRi+MDR5k5sddxilwzpZSqCJ3WwkmV3O3X+eSWfm8GXPpnEg6re9I9q
W/Isb3HdKcy+eBd/Pc3A+HEiZY/ZRZgMGgETCLUVuDyBa+4eDRbf8ar9f9RksS3U
p2xWkUGKaVXjB05yZYmU4gonTDsRUFd/qzemnYsIKekyjDdteSQWVyocmPh/+/iz
+iBVTxsAoUKzhJ4u5ougFp5o1sQKj1fqX1whFUULEQG9G9ViG97hVBUhCU40fA2B
K8yFsJOuobw750hwNmnu5oMVZuywSHKe76RJZqIGbkhYo9+eAGBH9RpmdyRRrfCm
B3mcJZk0/bjBvsAA1EGTsEDet15uatzSIUBoZhemUZ5WFDREgczdKK/T9McEaBfM
WEDWnrF8q37DAFaJV3KbIct/RatyjF1Z0iDRrtaaFvhNnaYErcw512KgpM1030iz
hkKDWvto6hHnV5hv76v8TWP1Os4asR4cm3TZsnHYen27iDcFarqNoSWTo0hIdkXe
8GaaQbb1KNnyjo9i5c9Hpgd0ZO0SdJbUWL4HGfzC3ABqs37VF88LEjNHN9PLpC96
2EbpJVi1h3mPVQDj1wkVb0r114KZ+D+uSCWdQr+vQbEGMETJK2pH//x9Cbm8eemu
UwhleSfQH8qcuS2aEO/4tVpHM0SVuZmmXFIsqj1gI9jr8LA4foxNEIhcot7qWI91
96IUnV2DIqUuusgflIgVPH6fkOMUKbJ04QE9BAGNPf3dLsR/xa19htTkSI8wPoix
iMxTg24NpF04p3jBRd5eqAplJ5KgBfdsLW5HnGVJdycnSfVLA3fVzumQ1frC0J9a
24/fxdTiY88gLG2BW/bQ+axejLLVj3OOPU5h9XPbLR4kf5cwLkbm5yH230yJnh91
ZmbQno37VyjYiGQcp7ejHZihCWNuOkAT7RzvTVnP305C9PLrV6zsxFZ9vKnmBLRa
CBCxTWa6RjNHMTpLhzGjXlvplvBJmfh4rjE6lsNcXX1TrOTrPCaAwLWKmj4iToFl
wVktXExnlddghXLnyeww7Q7B8LsmfejxOJtddDBCCyfNn2/RGyjwYzNnXdsNbQfo
UPb9EGJTY8//qBe4hcNwYopQvE/KjAMu5tjCKU2Gxh5/Um5Hx5fCOSMXbxNCtVJq
Qw/Bhj8XNH3AqOyOG7yXfd3s+68wR+UQDc0aNlagugFbQZ+hSAv6+b++TKE1fzun
Srj1BSxbEw0T1tGMYM3uI2v/NWaAQmdaM0Zq0TEtU5Y7OFe1IEFnhNsBSE1ZA6U3
MBYPmiGIsHSokP1DBdJSU5pbXRirie4Y2Lz23RBOys9h/4Hif4jcYP/7aINf+ZLJ
pFfOmF/BlFpObmqZN+lbOL8MIGyvWvsVGuyna5Px+n5wcjhe8YdzyyRkBetDRtGZ
jpPe7xQSzLI4vyREA+ReEAWLHXewZOsmds+MKSHLPhtqHTbh4LwGLscbmGnA4DYf
M+Pri9kLT6TLTWDO3sWyU04bvCN07bbWRmujVQnRS/Zwy21swKiivPmHMBizPbgm
K+JkOqRTyRQOrBtqlrlwC9538k2mkAcSQdausG9I5Hub63u0k95fTCrRGVO+FMV1
bsZOUL+HNol60CJRFHVgUjxsE7AVOkaedh81JKoPYDH4V/tTA+uCkigkw8VrKAzD
ef0x+Om6dsVWD24ya8woMTzNDdPeR3iT4cyLh/5pLOJlok69fXz/HvR2tIlTA+F5
XGcZzmIc2n2QlzKoSzhVH0/fiTlCaRC3tY2FF6PkiZjQgDcITPdmgMsqWZ/SSpgs
FZO6CL/bsIRg+z7wA9ACmiFLMVn0NrFUOGTg7Z7sQC5uauF9P7YjoydD3wDUJHP/
ltHuXAaoExoojS65S5mDc04A7ByW8ECuZEeFHjbe5aXPJGyO+23R4f5/HV1fX4Oq
HdgqI6IMCT+tm39IWSD8yUWZHUux/IIXWZ3sFwbiUggkMjr6AIkyHFdHjspJKJxz
R+UD6gb/sdqiEMapt8PHt+8DQO4OoHlLHKlNfzz9eSmBMwus4RoAmxjweRKaySdI
e2nf0A13F+HZ8bT2SITqsy3NcIXdnYNPJnREbUNsp10s00KE3ohTJKYrhJuuLDcx
AIv6t6OnXpC9CPDxU8z0bXGx9wxWd58K/drOEmfC58QE3VZOZP/JiPsESqZ6SBIJ
wamLPJ7h5iirQ8DnIwTbDYXkui0pDWn8peRg9xkzFXYlSNyhIw0m2SsG2IvuwW+i
6BAzlLQYAo1C7CnoGzVxf7MasKi52H6IBE5Ht7c2Qp0kuVKgvlCS4774qhNnuKez
9bv7PgwwkM8qFfywl2llPSLGWT7stBrrsq+UHdCNBtKHk7GVaJ2Jjk8B+ZjiAU0n
DCGDl/m/TDko1WE9nXWF45hV0RYAwrmcWN8oLG9CCdlGLIObImE681aZXQsMzchc
hywfsfRuhpyUQ7s6IJVflI/IRFl3ag72AzNsBQAiXJrxPYwti4HFVapvD4/ciEP5
MZx2KfUuQpOngB5iueFVYbvrCJZUuwlXA4INLsMNar83R+ex3a2KkgyaF4C4DDW+
TrKrllOF6INvBDunexjvfh0xIEq0Ug/vUzKMfRCCl/JtGLuzzRWbOxCqM8PYF9LN
ymZFVZSd/OagyMQnUmATN6Zo8yOgg6Fcx86TCVR1L7tFiYJWcHgNpydWZmBUtafy
yfyNWrK9dzF3zgMGVdv6xAFCzzVaKUaBfmiGuCLg/pwMJ8YsMUs4SY6uK2vA1un4
QDkRsZH0udjE16uVtJuvcwSCe7v79UbLczBi71n3BqgsOZ9H79UdaNV8b2xLz5iR
F0QALpiDyOLCzCWd8hiIm11sj57g6WUhfh7Up1kZMuySFXR0Gl64e7q9Rb+w+fg5
CztZ1ZEbRMHMxHGiXGq6ZPLhZcGg6+tHBx5ZGZIFj+lSfjXyi026av9diqXptnUS
OFWiww4/hLzZIi2H9yfp+8claf7UWbVv3LrnQcQ0Dd/Ya49zF309koSPJf6pLAmH
/OZvyAffmKY9WR9YQ6emKoLKIJMYGbx0UssnLwltQzLHvY0X5Rg+tKCD3di31Ut3
aZIZ+0puSciTPFdUuEgeHHosgO2YeeoTMevUDvkH1I/ehAg4nAttw8tKdN6s0rog
PsYEN7Cnm1tVZrdMC+A+YCnWyYD4dAErFK554u292XU0KclJsn47g9VbeTBRdKye
Ib2/izRUANEMn1e5r5jR4OeX3a0GIeelZt3UfuBtKwxtOr9EG9L7TSrzPQtfAwde
uJPetE9yMZBe9XzGNFFbJw8hCzwjyOAlczbqp7UBG/BAvvVu0pfIY5TRoiERT9On
1OUgQfCF7kAngp0yNuxvwlSRkFJ0VtSMP6kv8whWxDzPflndBtI25MSOqktTmxkB
zKo1kQATfPuqW4I/BTVoOplTICCm50qnEfw4YeTWWuzHB9e82KTiMbrNZxUAJRHO
8b0ndqbYt2x+ceTm86Rp3/ETHP/DSOtk4gHxmsFthgMmnQ0e4kdmCCbgpbAdVql0
ZTFKy1LcNs3Xqyp1TUbyORAEzrtkJaV/KwOk8oDwbXBhpOwYpgrl7vq+fjq5QzkV
2YrwbwiCtI8X7pkQJn2DKmCXNeon/wvP/nXqD+caHGkzzDQ79CweAhCtxGVM2jZT
5sqKRG/MOWGe0vdYVtzPmYzx2SC+1b5vPAkDUbyro4SelnhSs1b/Ghzml23fF4WY
3qUcxtgde1SF6Bm7QBrumNaNwIEiT/GiLfxp5GIDgeN9Z2YqbgTa0kMj3MBZ0Q0D
appEET9kvmHL/Dq1a2dfNqcXvE7vj2mCkBO5hXzGK2EberSTRZxzW9GHHkx6nE0h
K6fMT15fh986Mr1GG+ZdaotTskoJ9yG8DuqgKA8+vq+YqoJd3veBGOYVwaOw3qxh
H9zNODR0trW+FHY1NodFsbEZUzJnYICEqGZoh24iErsLGO0zaTj05lalSVdxLYG2
SL7a4toYpFzZF5LLjBKQHIOgKiXPMGpce7oaCfijoIZ64x+/XgBjx5ddRpnGQTNr
KfMaWA35QmEcy9y7SZUlqe3EFuG30yYvN+yXSTD0tP1aqlz1e8z3lFv9I1Ez6Xhy
IBdvzLCysi4FMV+PeSHaw9weTJ4i0vFalom20o665GE4MEqlXZqpFok4MDi0yWhf
K3BSO0CoXjqEmZSZZ3ZElfaVMlLqmeg9MWislQ1Mp8duLop+aCWyiJe3P0gDEFff
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
To7TAPn1kF4xIdsUS9NsgzS2M4b1HPgq+YRKoDiWyH8ScuZXitYBNvjHI8Whemxk
1rl8K2wzzT2oKbXhEWaiIMKdJ7lSMcKziCKFw2sUHw2uLFjPDeQ+2G5mtbN4jMXt
e2CYz9T7WxeIGa/uuhKFVQhY29UqlakiAdh24/GLaeseRbN9fJkKYVgSj5xObSPc
aqwpa7WPcGbIL3xGVTQ2G1Oqjqd78qiV2kyo5VRKFonT/otzFeHD/xluL3WqjYPI
+FHHPYgo91793jV4Xp1i1lsCTXxqRWKGQtal6STFHdAsK4iGUcVZeN9OcyDRFJYK
UWe1RTg5PRJN6AEwneTplQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20320 )
`pragma protect data_block
Z5OAPCB0hCWSbz6y0hTHx3CAopW3UDIPGX6J2m74VL4drcGMNNNZgCJ2lugXErpr
7otwcUL1SjGKFBYGHiH6m0r7jxEK7w7Tcw93AHF08KQM6TNZ0A8U+yFElIeWn73x
ewbF+oRZrqvYo155OjcrR3TVTfxp5idfLM4wC6xNGopgfPHS35uMGOvol9GK9NhF
H0ArLsGwZRZE5iK+swdWf+edKgceFlYIKpDOKGLAfoq+Nh9YxUsjHtNK0wVtHL1+
7RLUL/md04FM/LlzYKuj0FpukUCHxe55rPkMpleJTQdZgvIMK7REMZrrhaT0AaZX
olPstWwkuI+G0xOwzRFAgjcspOUn2WrJca54lX/LUdys8HE5HcAe5rTeV3jTIkCD
UUgfhg56PWtWGPsP9HqauLi47dayiiIzAi3FJhAeH6js77WrkYq6d2OQP3sgiWM7
DlxtfTdi57rVhUVrSRAMUdg4HpVxIBYNxmWbJG7YD9JvwkzItuulhredJyR1eM4N
8pyrvTHVpaHlkpbdzMQeXEZ2FHiyi8hSAN+T0gOEeub8Kz/POUJ7xxiw2atDxB4d
8TQPbw9Mapfa4o/9I+JLBHHCscBUmIJgvP7t6w3/HZxHBOskg5oMW/JV/pjjxNDs
UntJFq8CsB3ADQ1JmhZNoLnzlutZBnDlgQVZ/ItfAhUpj7i5n5duWV0+CMCnKIt5
xoIaVfTECnYSUhFTtRb2bvw3cAhRnZqznhh9XkLyGHCeITnLXuBAfAohkV8hF4kd
vtDH+gXSn4Ey9yxhYmDsn1mpQyxYCikwosQLJ71gocDiPU1Lht/C1qjZfpKNo4bv
CckniX2Ur2Hs7JGN0rB+p0GTnmg2iDh7+puHUyi8P57QS0cou3TlxfOjBXMlZwca
Xgphwu8fbFhUkc8R2TkcuHn0wlMuraxqm1uwn7KlM3Mcz7OoSK4QR2utRB/Hg7UB
00QBk8FZyxmLREIpVZSe14GL/Y9R2cfy5l3OZLbPCyfjWQ2rLaXMeazHXv8P2MtO
WVJriu4OdnaLMJOo/m83uPkECl9XqNaiM0cId405ANTXpILC2MgsQ1Ua5L/tUens
/IIjP8QgW2voFo7pciPDZAgxQmsrUoweX4LumTFfNP+9wHVTSQcXqZ5GG9urPVzs
Dgh0WZbgI7YvrQZVXo6vWjTjsqufsVeVr7D107oMWFQUUDkRLt6zvVfhhlXB2pQ5
miQCkfiSG+HGypPDJrBfucSjlpqXK9ugrrt63H21gVnmTNK21h/robxN8ZulyNWC
+yurvXzvo5EQAShNEgeHE1Bc75R5D0Owhgwtfm7GEAp+/wOigvfx4kwNm+0VlNXL
epCT1axtot8nw2s2SZHWe9foFrirjBwPiDU4IFCwSV7PlJxWhVgtmURjuw1oqBh9
HdxYjDPcmPK4eSzSCdU4f+xVa5oCAFBGdTtiJ3/tvVs39cITuNgWGMZd8UE3HDv8
xsrvDhLi7BeYcSlwVgkoUlN8s8Txxxj5lG8BMB3BOINidL69/BMZsDiRPHinHnUh
8d6s9FNO71nl1TRLB+6Ra7ZREN+n1JhsmY5vGe/ylpJrlEMWwfdfv45LXxZIc/5a
B04vgjYJWmPEfGhqw+V8bfiOaRUz8jWioXBj3Ays3GZKEZH8T9rxWGrLFihi3SAo
VuVnI9LS6ywXdpeav7gnl8bGxIQPUD2oxmJjiWE7Y8ZecksmNgMqUqlgatBogjcc
pJB2az5yLGDyuXxScHycyDiLt7AAlnlusBvKYFGD+8Xrei0cjogPEVd7kTFtWiSO
L0il3L770AuogxTX5pZOcre1YuhcvAMzL3AQf/m2LAjFLKxhrXLajuqf+0ik4P4k
L+sRJYVDHr173AKn58BQ58gOxyhK7R2MFj45U32CAKFGilKBwO5XlyURv39moJ7N
v5+2ddUVy37+iouAv20/wj8x5wE7KQKw1klydSyRShbla3qSRiCNr1qnYufMlPIk
uVtqT3v6P//MlD4iZxV8II9JwhPo6Lju8w/D+wuoFWUrmN9aHag8J2U+WmzKONKN
vD/4BURlxqCjHC/TsqrxQBnlcRCkKIRQcNGDLVo1WNPgXqdj+6UlR38Snff+evdR
Jk0ZtL2jONFW78nTmxp34prUcdGDecz1nZJ81gygXoAN4fP1FfVWJraZoQ3ZG3xJ
iinQu52AAVF60oyxl1x8Nk1aj+KDtRZw7sXncp78JECOxVJHOrUdtl9TfZW1V4RC
h9ZFnHhuftoq7q6JDMmJG20jTl1KgiqnduEEHr9du9u0qw9BN9Jc1AF6fF2Cbhhv
a8kLn9/Evra7buuXlSRyOauYm6MgiIdwgiVFGBUiKFaLjqOWIGULgzZeKoD/X0pv
wYDy2F83jA1IRoqCztgPitANwEK0XVhAsg892II6nyik4TOeGjmPrlw9C72JPCX8
NfhBLhLUr9jsZr8mVpYRfOXWMYUs5F+9BMEAFKvJDX3xZSJ4s6DiJlcP3aDI/CLd
KerFHQDfI4sjhokzwyE5WoahJjmrZ8tcJU27ll1Mtp6XIjw5ACmXiKVORsmt+qzv
izquC5b666zh8RDLkexEnVL0AMnfWKWxi0dkuiVCn7c52RaY3N6XLSLQiU0s+KYz
NpDVvtRth87qx+77koBpfzOb2F50sPjZ/BnqiwpoO8kzXyf8T6yDYhHKXueqiWOF
XvbwYzeFkHQNY2l6Uk9/QMmf3MQ2Ed2NWuXynX0g4UtAs8PEc3JBkDlS4kQZxUOe
b5su9/V4gizrsv2rLOHdolCwguLFg4Z9ltvI+067bBK4AFITAaN1iDfbyuQFH5ON
TVhrOiNUToN+GYoFNPuQPnVBa8nt8x8HlLumXVC4nFR8/AGekEXcS9IW3Y47jDuC
EtVomNqzsiXWefDLJsnji33ZA3QL8OkHRpIsxKpviqF3qrOviVkGwrlfoJOGmm+5
ficHWCCfwzaJ3Bwih20eOfWxq8JvwBFC0cqyVrQO0l4lYhP3KEwUIeVjAlNWEdzb
WYLmemH28hVeSbcWO3Zz5s4aTH1nj+5D27gmKpe01u86mRlnhQblLfeVn6YnhOjB
r/uVeXbVvsI9g8RmzNPzQVTyJWrqjXcfrB+nGUarhkccMsiu+5QLo6JJlSH6fmkC
Vzq80r9qRFykKpXp1wl750/LvRtTIisRBgpuCYmdknRIMr7VdFGMnZTsqA7NY/lY
filTl6j4ilAkZ2mXJGS9Oj8Ih38TSaKKMBG1bVrFwdjn54HhwswqFffBh/Qe4ttf
0xzLvOEw+jaWQqataKaq2+50iEQq/T8TwqYyY5yzEtXtPVh1K1PyjeM82QszAS6Y
bqnRZBofaNmluRDFvB09CZyKcVXdSH76CtRZT+QYXNQBby1wYC9bCO/Qu8TawGOR
w8T/iNNM1qqV8AQJpSGV8D5d5WbluBCSOTyLDion7oFKUZsi/4UwgvAM3zpLTYFG
UANfd+YS8nQQ6jVyS8y7t07Je69XqubZK9kfhpcxsN9c4iF22B2meua3GnXFke61
In1KJkXPSnJ8gGYLmS4San4r1GrrBnvdHWrkWEKCj6uPuTnfGh3fLluWpf4hBN9K
uiyWIZfeUZZePuHnXyXFZ1rNIAW1JY/s6MhEjnypY0WIvqxwZ5jmYXN2aT9aOFmk
sxVjuUBUORjWHZrjIzf6LkwZzrjq6qn/YqAAfjVhqFfHxhffuwqcFbd/4uleH8zP
ktwXDLnn6fn9BNmmzePAcUZKppju1roRq4Fg3WwQ2UTMJTamTBKnEGVfYiZN+iQF
EHtbNNUZW8H7xwwL6h9F9MMC+FXs8ppTYZDOiLNfHzrjQ9tqEWVpkiw/JGE/QVm4
Z6DMcqNCP1xqhCSgjJqo/idDcFtZCCXsGpmJXbn5HNd4q81BWW3StaITDq7PF7dw
aqh7G7KnL40Ry6SPnWewras6Mm9Xoo2C++e/IBOhy4QsT9qOUGCX/7QNM+l4Zq5G
d5KanDwz90l4q7FlaiqQCLDGVln9b+s8vd9AOIoLZlUlvJfbv2gJtNXLsRWtBexU
VQTJmxZ4Xp9r5ifsDZ2Rogmc4n0MNywk7fM/36P0rwaE/UvJ+Rna1ZCy3iVY+xIN
DNzViYDQqQfh/vexs4pkPrjzWT+hVe+cf8Mh63A/SAkUvrWjOd1l+CaC1jT1sdY5
a5vs1OoDKYdtAGcqh/Kwdr/30nJWBA3WXw1UX7TWosRIUA5khWnzuK6vCvhPbbS0
NMtL820xcpxJyV7FGeXFo72o4S2fLzSXO104TVPE6vlHWl/X473d5hlxPh4225T/
cwqiDKtkU+JhpNsN5b48eaQGqYJBTCiGvAVEIRIsBgPddG5bx2hoozlqZnNvNPzd
I8+9BvVsxOSajSq8LC4Tn3R0FxlntfrVdC6F9QaP19HWZhUbjeN0Bqj41iSVCrO2
yLsKlZNkh8jtRc80NQrZNdBNzNyDTr/XbGNbob8COIymv40nnc7v0ke7+KjsJaIW
T9AmmHYErOll7/kVpt+Hn+5VZJ+kkxgRNbvtYd731jyH1XH2uvDZPRwfjC+daLOi
MXeXRVZOTBeE6qq/i5FwZ7pm2UFe6721J6AIApNp8SGmYjqAmhuu6SVSK6eZBTGj
TQnEI7eYB4gCBjMTC3SyTMP1LDNH9IRzq7eAbefVvCD82fDMYuCkqrD2YVy5iix6
4koIrn6oJrP4YKChvzTeSZykxJf0oSRCbcXPPbIRdWXqXIE8MxywOZZXO6uoGlJb
cNnXt5DtFhD/ytt9JIO9kg6E08JNmKIwDxsFEewVNp0EZDbWsEyx8hUMA/SNDnj+
Z0jcAC3DQVp4zjWl9uXCofO/cKxX9vDEzq0efY/C1QwCjvc1pE8H5MHTPDey69+t
8MkbU45W+7sfu7GAVWC7seLymF5rWiQcxHi6n3EPxQgtcNKqewlrSNfw+wPMsRl3
aCU1dDLLPmXH/F9/Cz0LWqxIpgW2gyOLdL7Qxgl4vhtl9ynFTA5HGCvu8yPau+zg
dxvR0xxry9epwW72QQc8Nh4paPvTZt5CxF3tADJYSwe3xri0K9rg+7IQaULK0LTi
xngVUC4x6WqwjiqnwB40pLDDvubjWa52mw66gH3zZgrywLSRBDujr0XPDv21jaup
z/vIIFMwJfBMj17BgF7yUwtwIfBLr1kURtw39kDBEUjPruq3R/g6tx7arU+6lMLA
8oDE2wBnCwj77Y+Ht20bB9+vMmM3bmm9fvoD1S1e5cESz666vegf6+JTyqc1cavi
2JsB2trfTPC6js51sYl5ZkbRWBGzfJG7z5dnwzXtDLmJjWw7z7VNJ4YLTIqDG+it
6WmA3f6DTodEGavd3DT0N+FTrWyCETUnXWol7Rf2fR6WJ4x54VQwxyeYCh404Hrt
cEylnkXmuTkWIeuSLp1O0mBGaYC9xIT+YEngVvl0Karq58Gi0yUOH29u0Apl/+bu
+UQdqz5TOVWcQc5Yc3DNHKwHX8v1GG+hyLwBPhVMM1m3PQsbLdYOlB9LNfnkKd9L
GJvHXL8EMkC7k0wBS8I/U1X/B5AcTZ+TVC4HgU7ADtKm8V35U79hRBU0ZTmShirC
E8OH2IXK5Gf7dZONLOghDLZbMVLdj5IoCWHse+XIXZQs3IzrgYXacmbCd4KZ8Cv7
dCQp70ti94d/4tMnP4WIl6aSXRVzxJFe2GYX7Ax89GLTfHciNKiNHlwVnY5NN5vb
ry9WC1IoJa3Z5beKMy9uVHK1UdmWYlspzkKX1uELWS4VzSnYey4WlUKZgb2cKeHf
0SVOjtCQBHQZeQRlezJJYm/U6w28S6XkaS+6UbG361liEzX9avLB+N9MJPyJledH
jgTycl4pknCHlom96lOkTjSEcv4DGvyBWzOi3eW9GZKCIjrB2Jvn3hg8Z1D+XcDq
HSEpqh8E1Qv8NyKcfOAuYzlxBCQE1F/3SPnDzONh7NHr/p47kjn46f0YMKc5Vcof
+DZRQWIqC7uCL1unwE0Cth7zHo8ksNpyHV3Uclu4cDWduiIEFuiXzPj/cd2VVwxJ
roQaoxguLpvAqJvGACt1PqqKeTuY5s3VH/9U0Sox/n/M87X1j5Rkv+H/VspVKfrz
4/e2NFrQdbReItuLO2t0w2eIC7Wfi8i1hEqUbMcsK8gHb7z+Vcu4O/Es+jcqWjVx
qKqBTUQ1J4f8h3IvLkyFiunRFLVNxpaiVFo3GIkRJcXpAohrfD07d3iOpHXbcUCm
2Xj35iAJqM6yqGG9R7UYoC+IFBc8RD1VeMOux9TJK1iNL3q0BHYnMlidyG/oo2Hv
ZCiSrbALD6RaXpZNkVNjIGZbE/uF7Yha1w1U2OF0KNdgzvEHLmbA55+tUsH8J+7o
rbVtzgaXtwO2yqJKwdZz+7FhJQJCkRLMDAQWJqOyNnXseGUJ027kOTILMForrxE6
rARBMEY8S2BEZaZTbsv8vGpMWo4FvZRMmX4kKm4gzq6nIeWKY2qG8OmWccEEThdo
hj1Lhm/orpvhn//TAgW+XHzjkpfMv/kQTkWZ4ZdlCxaWhozw/guipavzaigiRl9A
OkzItaheHHcLj0UwYLHtQTm21ZZj7Q2Zq0uvAfiDui/LgUgsrgznKhNWeqs7pyRn
D+xXYIYtKgkJBNgF4hlETADsgOQVlJ4WaPqDupUFN4kvcL53w/fsJrGNs16EVRnL
ukCXkVequ8rObuR09GnECQTK2bm3MGqPO09evEJ9pGTd1ovprkReWmyBjGjfIbnH
xzM9PrbOVs3M+ENiDC+aRSBQbjhkFDPLySofmwx1G5U3GShv0RX0mXZGadgiZtn1
cZXxKTWkVyW2B1ywr3FWa8fsGLviskxuJnNdXW8H90y3gaQ1NNnn4g/FCo9s1a4P
hA406c7bhG7zjIJE+zkBWfTjjoTD+t2zCiEXkvJJXApF231t2QhIuAUL/elMTOvY
CpyxjKCKN+KsUOr/FiI3OQgG2DmuFhlCjQOZcdSpExzLnfTw8PdF1m0lCcvz105H
D+CoFO0EKFm9bzYNO10zm+qI5+v1+C2vJn3+9e7lNwNleJRFNYMtd4dJ6bSToggv
dSA0msdLskUrhm89xmXkY+tDNN7yQ8U5D1yMVg8HYK2z+isTWOsBrGqZzSTOBAlp
L3S+pGWUL3MHzBxTyvK8a2O/LFd6KcQ1bhvCaBdNhCBCasSahpfPlGkWGJi8qXX6
8j2h/01FKbMSUe1rraPMX9JlmHv/dtFNJEa1teRNvz9826ASP1GnivMwmjH0MmnP
bR1Dvdt+u00ffScIPg/jKDKoCMq+/hunlUk9aLgKf0SmlBLnIvi+/LbqofXXtKkD
hUw3pEEIZ++PPdRaXYjIoGIZHVrmJpD+R5BlQDdJX0dbheUnXyD3DBWzf+eegS0r
CltgmetSB0skXavPJOzqMu/eI31P9K0weK2S6XPJi8k8qnxZXW8BzKkldZkNpf/J
/skVQQeDSWPNewpahjAJGNw6VnMP0M+jOdcseXd8FAfR2NXCnB5J+mvN3oqNO1lh
rVwEv41eTDzxs/YqTe5cHoABPeLn9Sw/LhtAtDyi0n41nSjxFTnT5IUNsNEPQLBt
z5uCMqNi1F0oSU7lGlDZuW0sKgN+gPNk+ByteYpSMWg2DXg08VNTmVLdljtAmNNO
lsT0jFFJJI6BNnuslB4DL+VACmU950MW5fZAptNl54lHbUEysCUdX9Msw6ZofW3V
n+4OJQGFnWXUry+JotlTrQ61osY2q3rsfnXfwwSP6gHSzInTeWmdQbbMTLmhqmW5
nH7U5F3dtuzwkIX/GMk3qmm1S+5w2I2iTSUPSZwXdx0+9QgTDmRSk8TAClGIInWs
bwVgHNxUBFJPbS07UC/30hLrTKBzdc8HTeDiVGos9EceGF6A1ykhO/xRFiOvMuxU
ibFAY3QpjKP8Yzt4Itp+U5X5hdedDZGTr4u8AIFrimAjhYX6lg4/LmBCMe+Ocd32
4E1DobQJhHXMFfhZ8aMFlaWtWiuBeu1rmaXTWZkpk4ZZi8RA14ZP4NAjXC93E8O+
lHLxs84zLUgWqScea4S+8gfaEqeKR61GDblFyEvP7On3edHMRtllJL90ZHg011V/
ftBwWO04tMvk7iHh4lrBmTHnfqSxGCowfufToJvMjpdp6s13ACDyKLq94meez04u
XoVUJIe7Q30mGN2Z5G802U3i8tthJQ2FMCJV2cfjPjzAkin1m5QUggUrwOXuu8W3
Lq1mG1XKiTsSZbucVMPM4e20DbpYVOvnhwAe1+ENGdt+DDLz8vwzPbqdujFC8WCr
dpJIM8P2W74A8moy/KLQEKJQVVcx+ztlPCcUs7OenE3jF++/RIXGac7HgwPxsO1m
jDTFpUcC8anEhTGAcp/FAGIXZyML+nhisBeDei4eqKXaZ4c1CGB66vmCcJ5IqA+J
0Ft3cfupxr3zvwZ8hhmuNxtaN7fVgzETtK9K9ME/NAKBPtMQVczlQPtYgVaHmp/P
JkrgV81QihW38LwmOmwKSBhBqUVLS3mpOk/rm2k7wKogcpaHEtYmu75bm26UbI3M
bjCW5DFqyMYepuHKC8or+oInYl/m3ana9cWOjqcdLRYrBU5cr8X2SQXJEGRuzQyU
cWU68qdr0Mw3ztXKAW0jL+NrKWI5d6mYFxzdw+GEEcsxDAaoaMd1m/bq2nGnBl9C
5NO2PdxBZkPse1m+ENEdG1LJB7xhDDkxjqHbbvZaaXbUwEeMJZnZcOcl4a4t5ufx
izEZbYoTzw3J0h+qyD/FxswuIdMRtTFQP6vxS6yOGZICVk/fjjjPNnMxjpBrI2aN
ChTSXygEymhIb5BpnegUvnito43WW9bMF3vwGqJfYQqDd4roSvy2kx35WcauJb7Y
/wNRyeU5bsXR4YGC1K72vp6AtXnF86laDSv+s/bi8FTbjIkHCNa5CfRkjZkZ0P/r
Xi7Dsh5+2uPqOeLAmEKzIfdfC/NN1Pau46F0jBrPQzURp7kiJcOz3TzSCYzf9dEj
AqllKii7gRIOcJgfWC4rUyhbIMeSFSxZXCD90VneJD+1N1G7c5RdY1k//BAVz3ZK
3SdNWbfjmz7ulzrZFVYE0OHSRvP4dt4/j9ETxjh0gkywhFXG/EeReEM0KVI5cUdu
+ZeFsMzKGDA5DehKBrphx9yAXemdNfst+073E4Q95JWKO7qpNmwCrJlezx1XXSv0
B/kLDMVmUa4oArc+uXHXLFBX1EGKCE/90DOT3fUQoeTiSp6IQULCWQHgZP+bhzP6
K/6DzOKwvaJMtpjqs4Yf7P9PRXy4N8fMbYm8xaJtRatxsp3NJq6f+aoZsDrRiysB
K+bxY3DlGkyrM4DnOHgp6SSD/0OxYI/I93bvdRsF31wRBx9f/iQ8ljx4XTeTEg4f
3SyVRrPqnAunlkEYTxkiOvdtpa68GQFCKaBWuSR6tVBf845DY2VO+dEPgnKqe8NK
4nFFtjbzsQpfG7aFEpUb3oC07F9i3jv4dvok2hVvRYDRPdD0EsVpx7LybRhAdPt+
rVWL9IhzS35wpYcZb1P9o5PC+8GIx7+llrX98FULwXamgxS3IClIn+3qoxeQr7d4
1oy4e6vPMt9P7BLt8fJ+TgIixS4EJjeG+SMXL07SDhrFCOWdrj4KU2rGkSkxLGeP
gKolcsRLW2DGvKmhbdHtJZJrIpnhzkD1L8SoQeNdCTP8X2BuxDKceGmHfN7JwMhV
rWPAfRTYOhM2v0uU7POTnQuc2/WlxBjo66JXWPe6XBDLm5wLq1AoS4OrqRIfXoNU
f3HXWA4bfVtr7Kw1vBCMgNAjV4lWv2K3/YayWWU+/qGMUBPFjsJio3fw1AWfEECQ
2x8y6i99Nxbg4HlxZHD/IIGhFF1eTcUtYoB8x0QnEm5VRqDWk5oseHcQCgxdMPOD
Pz8NueQwpoyUKQtZM7XRRh8OcH92TaZB53Mjzn4xNNgFbjjzOQ8XVU8blSVUWe+E
SLujlBMfl55/gNT7Pj3uucYGlGp/mkpS3S7DfzQ5ktcN70tScx4KfTAwP06K6qlz
0yfSh0fym2vI9ky0dFk1HgtZ+E2LKncTEjw0npu7j4YMg0lmsREdgehFFZIbZ04e
k4MuvMv2FlqwSUvIfESeJMJhX4C+gs4jW7yLpzGeqz9TyIi0mdy9sQqizqtqUAm4
NodzhxGFfEcC9LJY+sBzRNA916M3KZiHSATVTjizNYPBE/etIUIidcR8NMf1xhOa
FWKF8FmwxuQ8YW/uGlvzVahnslW/CS/IrO8rS0wz4NGtU5rVMLejrCCNGKhKcJnq
2rE2Lm1bX9U6kpnUZfqkAuTXnalqzOOFZUyLItasVUsaolc8HZPPTnJdWqzoOnee
kO7YlufYmS1wnuH7FufwukOGsAQHYVa4eOlZ4KQwdZjyP+4HhwoTTv7jBGD66pTZ
hreCdD9V0cwZpzE5hL27C2xpx4zJBBfrdBTbeuNZ8cNmQMViplraN2461GAb5yvp
W21TCm42vk1xSKImVJQopHHDUU86zj1LrcdP9DwC/iVfqdeyuKVjW1Bw7C8cRn4r
t52woXBF1liah8niuJyeUrDMBcXotVeXHTPpkk3Swzw0XmTcnxFIJXns4gd3ks6/
Z14ZPapbUh4lZxzSaFvjvXZfTmjQK9trwbkOcx5yPnP+8R9jo1/cSkogV3Dufs5D
Bj04omrytBrPoePaF9PtUo7QoF+OmsNNFjHL0TTwdBAwh8CW9fbTgnjoJR8fo7IR
JdSzxYHdwD11APjKc0PvqXVeutnPkYfiEh1DtI8W8MY0ku2W/WodMv2kRk4QCs9F
2S+uE1uKcNZf2XL922HN0sZ2Lok5PdBHBRACgv17aK4VStljDBkdtBEK3FfU3VaU
mvl+USNmND1KwV3zi6dxZGKhGvKDqegqSiv9/LvtUvKPLUNJcvxcLjl5lAk1WKp5
tS6B9J+5w4CKJVSXLGvb6R8vUcV0VAuHJB9+oNIqg+sMDaz9JVniXGQdPX2ZG7mN
NwcgitXcMU70EDzyHitFYD9lutwtPf7xvpX+j4lgNxZpaef52sMwZoBe00lZTn7C
j9sEX0BVxDRmLSR387JEx8ECEy9AXBmwW+v5Ovampzp6RnOjvyGMgw+Q+F7rtqEV
b5xdAnQVhnqbWJ4YyL9zn4QRSZCPWYmC0NFgnMqekmZmse+xD8dJhp1OAqAekh2T
ajht8e8+N4crlNycDgAaEqpLWJlpfa38dBwtW9VTKILV+yT637LQHQetNeFnRgcP
U6AO1HjPmS8Hia7WkRK39OgEDm8DqQ3neQ9kic6OtOJn5Jna9RP034e07X+Jl5m3
5bQUQaPPNU3R8pAUxRj0sLN06o1VCkN+bcpwbkV0VkOOPg1kOyMdONdSi1RNtr/E
zEqH7FFziUwpVynv/zhFU3Qbs2QOWVixh55pqyw5S2VHiAhdz5BxjOQPCFk7E2g4
J4dxTMG/4DTm/rvlmLlbuIjOn2D3y9Qzpy7XbSMiZ+Tj4YPuuS2Z1FA8YTrdBHeV
SWP2dY8ufF33Ra0Db4Ev+kDvsgk74soRXVT6595L8LLn1Dkndh2upqyqPJlNYMGy
Xk6BR4n7uVFwUvAHojUR2Jg8ZT9NWOlIBHOmIN0h44VgtibzWDHhU4lAt3ueai7f
9SuOfJqsNjFXNxFEtQEF+nAA+zq0Dj5+SaOf1O6Zg1Tnh63yt1MdlVSE23rbd6UD
Xvp9MW0JuFMahrGRLyHwBzQYvDevMXmbaGTZj/yV2ja/QzJVD1e2g8DIjc6DA2Se
lKaONXM13A1vhCz7DokbBeqvqEbS+YDmuGFdLcFCrlwLRUJPFc3Q+7J6uwo+BKLE
hRLBuUV6Jtwa3wPbifof6vi0pcytfWleWLGC5DJDxaaOPeyiztIVRq5SuUYjIy/k
pUTi4F5nCfRg5kbxcUxM1cYlQBt95aimFVX95/aaluKRrSEqeFe4dAIeWA9ZO7G/
kLKXyaBo44Vqw+ZTwGjfgBEFIMx3cPhCzQS4Oip9temiNmsc+YuCYDQG3o7T6qL4
cf3fU4SPQAENAjVr+ZWC6SgJKF3KYkmtSbRDPKdR9K3uHRKTiChoU5tHi0fyIJQK
OofcWHPwplYKQFXfzQpZeGvZNHq+Xuu7Lu2em1452qCtTgp77dJQ2udflnK8VhkV
ToRHej3m320f/n51vv45z7hbxGbwZBWrnqP02a+a80ZFY47NzR8ijn6MZ48PXRaE
8s4RCHgDDfq1dLIM7mJ8DXYrvYL9IZejQvbwpIRcvCtO07uNZ0cNQCdZs0pmmWRZ
wSvjl6I0dVj79bvvEFegyV5tNt4JSDJhnupXJcYRlyNRcn5pV7oiyiAifIJSCvHG
nxvb5raWATQV0e2wTT2V+HOn4Ow89xahjIxmwUvzwwOHBy8cPqX4XjU7tqEeuG7N
wFFrC1JVag/DcVt/vZJDrTza+vS3TUOPG48tAnxM0ycRxjO6WrK0hXktIeCXcKWH
jbqy5tzIyX02Br03T3A/yvU+6jVl/gJXXA20+Lb+M9Jb/+A6fGbtfAbpqAU3KL1O
FIaap04xN95l/dzuV99MI9PSdYoi6LhTciHG/4CVt87z/e9IRsYQLce+y2Yxuks0
FmFJZCg7HxGjK7M4GyoDfD/ZAlVf11vCdb7g0U4PdF4/UOf76odkv+WYxdV8N8KJ
Dl2Err6LikxM5bpLihwlIg7bjAtJGwFYAmDBv+qX3owhp+XMFgQcitSFfJQw4bXq
QutZh8exE/bVbmriJr9wJu6jnhp6j2InNGo7Zj8z2nvb479lVhHpaAvX+KBvYPrY
7FdpTpRcdWILeRHTfopAZv97axiu6MM49P+GftFlJyddsUazlO81ivmblMXqpPUL
uQnTA5ANukCw3Ax4xgQnT/uIJz/hjJ0tqwcVz2s42Un8xa+mboqCe/usnD7ey1rH
egWZAW+/GM6JCXjaTeqxCeUlrKy3jbgLWizeU8r+UE5/DYjgidE4SDLlgrLRXM/u
YdvJdqmrx4gmM+hpjrjYGmdWnIc20k31uFSGYnK7N+twCu9V8may51y+XweTsh3D
gcYgg0xhEha8DGmu+5cJ3oj8J8o234nhXK/DD84RfN6JnP01SL/B2psE9tx/mnR2
bCWFzB9Md3TsqlpOymYWFK6X9A2Qtlbc7LY5sERVO+xO2kdkNOijHe18IMLwZq9M
MycmuQIev+M7vID9qRmfnvwVIoMjLCrP4Bo+dT9ASUll+yFkyH07JxiwbtvfjrhC
uKHB+I9/NTYxqzQO+9C08nRXS0eWtpBYyLqiq5umuLo2vPDR3LEr7Jrljd2sewSe
kAwgEjbfKMcPB5nY2NcJfqIJMIrY2IPKDpgH0nrRty5K5o2TLTpa1GsK5xUT/ze2
zM2aQ8DamRSrbmET+3n2SnhArOBfHEiIohlzaF6oZUjZIOsydXS+eyfT6PJlBIcJ
1KTFu0M1Ty6QZXx+02m8mOBaXEY56HdN+EtZw0f+L+WkFEVJ7/Q72wp/x3nMV5yd
8Spo/2cNbzN6GSFBGqd1fc6twSGWi6+SsgA9mmK7uwMdoPMtsMf9PfYAzFwvPESX
b2lezJ0UK8xiQd7mtZ85kogmVSh3j7rMA/NEpB/7kNSnkZBwskOjEpBcXvBHFUNQ
lODRXjSLsnWeZdlZJ8G4MBgFMG820WLy8t4/n0L3IR6Yl2D8WaSBqoyrcxSCf5Kr
VRta6fGLEIVk2Sf0vImkCoLx9MEfGZjV/cSRIFsTQaORckZtId2uNcKdweKgF+rL
AiYLtYV4i4Ps2pmVLQHsDoHwQGQxmfFi9I+dYhXLB5Vy/2/bX1FHXQomyhjKankR
KfQaH9TtOs0flauHakG/QstKW2eMtkJ8LVIHDu8YqFMrRppxfQLotQyot7Xc3Ebl
TDHWk534iN+0O6zp0vZyr647iPq0WPQUO6JzhcB0CQ8VZt544/MvcBB6BF1nmVG5
FgPvUYjXTWQ9zGa8MDnZMKGdOwtGS+EKgOfDlkVEj164WiPKl3cS1AqaP/vNUcKo
FlyKAGPqXWo1/bA02nOeUAx2HV8aO07mH0wOBdakPJNnwtC3Usyx75zWEGRbmTad
LbegbGWR3wEarm+4pnEM+438MkIhHu9+u+XKZ4tXSeCeTVkDPEJ5i+6tWDzvHUPz
IQK5GrhJWsT8sbK9ogn360iD3ZvicfJI+RkQ3/5IFRSPhIfB4tKgXM66ipHcudj7
adW/HC88yQuhYCfUQU1m7IE6XkFXLQtYno38z2MN+FsuZJ5zPNrCiMtmi0hWMKZf
gNuw+kkL6ry31oBBWqCiKqhiincmel0wxwKQhpFQpWCnN9LHFnUSTtjRW4LmjUlD
F3qrDOLyopBi1+S6fd3vQ+RFcRWp+ZjhexerNcHM0d4yk/E9+yf5RfgVdKY0zjzy
mjKK6u5jMWMFLbjkmTbK29dJdd/AOe2LAtwbFPmruIKZsaYM+4XCEwGDIAM+n4lb
K1f8DF+gnOjF7bCjHcM4UGxS7WVyHgBQUo6DhG/Lp9lUOYzwOm7T4c8elxt7vBJt
qU62GAejyKL7Esp4z607KBUsylNfqUlPmUmalbhARLDGSjK5ktPSqLx15CeMM+ig
RaYU4b8zRU/2MZsqL9Yq1RcqBCRbCw7aqMI0BVjzfXdRlm0LguEvGeyWDudP9lXz
IIh9HidRd8Yh59KKrDsHHJmPMIGXWbkEqaZCDcuRc7mflOLCG1NBW17EluXkvkds
mpPcag4e56Zf3Ix0M2Bubmbbpg12ekDUrhPCnL+52KBiJ417e6BynRqPWUC5K/q6
uDQxvKkf8WnBWsrocuu1QiOqs4z+dR/AgmquohlI0iXakq+T4uip9RlAIrp1FZyG
3+/yIvAHhlGZob7hCiIsuc9op+2tLcE/GDeHSUKOUZ+5HRBaSQTI1RpTngBJt3gZ
HwEbhKZ1p02QEGKatYXU3t1sz84G/sQBYxMZJIcOaTPcemIfKuLKiT4BMQhUwX+O
MD1D0S+4Buj0mk/O+/b20Y5g8W65DhBuEzO1UoQAEzjaVId68Z2P1bxSEUI183Zu
E0bQx/33mo6IBxSZ01ehkBVa4GKbcbrUy4xrtyvgEuoAA3jUyg1gJGB9C4RfeSc/
4H6Uvo2y0cFZwLTqycJ6c0SyEKXwf5GX70cgm5Vx0rCW3tFhIQ4/Q4BxTzKzrPrK
CCE+Bcsg2m06D2ObxJzuUoPJfWlpl8bqhSLdM2gOc0AuA8lmoUTZA6e/+2HKxGiH
7mH2OHLTcuC9y6P8OqlqWZaqRxmh/7WqByeprwgUOAGEq06cpndfYQubtaIr990V
hTCkwzF80WE4DR9ziTFqrCYGdC8A7XIOsi63kkRuBJu1gsh1qw8ABiFTwjTRsGkT
1SeKFPHS67XCKskNaKPVvm0P0qfoI5Hyv4Bc8wOf+5JqIT8UN6cIfhkpnJDp5jy+
d3Y+oDx+4+/nqpuEWe/hu3Yj8h2+DokRha7PfXyx+nzbz3oRwJXFieVcy6Of1LTb
BDk5U/IQoYXBp7iax4GpTnhEfWtCLZMzEYw9thQdwPykCJ5XoUpAHRbNE/q5eIy5
Yd3qA8WstrepGRdrsBHG9RQse7YF8TxWFo89LvYWU1jJ5VpB2C4m3ljIOpNyCgT/
6u83NA1ESpyh07wYHvZ/PyiNDBnPY8tM5YZYSNTtWFqPVLRJ6T72vltkEvo0YCiZ
41XQELUEZcu+PWNSuq1tR3IkwJ6DBaFDDcmHupwijzC4jKh83V50lcgz+YhpOppZ
RiIyfYxtgk1PxgFZ0EFIXznN6RG5lBRTc12mR+iyBHXyG2gzrQStLu/cB8RVLXHP
hkMOAaxY6xpzZRIgU/UHA3hKg7RtcWq/FFux+nbvBvULMWl/bHkc7PBZidCTf5A1
F36u+BrdD0/uq4p4oSM9dglgvlCEmpbh84LusQ+zEh2JAMeekFyiGHSS+D+cBPaE
dVXQ6qalqtHhdzSXnmLIW5uGsu4Vxmww8gGkj0N+CyieJu38TuFVQafa/rFvm6JP
gXIbr/labXYlX4rc+QWJ0oXOEBiVlxL4QnoRwt5cOh0dlbphn3RprRQizWQRr+aV
4qCJaa+Ji6PU2T7UEwJOFraPxEvREQqwkN5k6qgu/biI9NsP7fOJCK7w+lbPqb6+
aWpXBdswbJ9DixAEuvlnzUZok5TLcwgi3rL+b/j7inZHBcHDinmv4xMk88RMixkW
tF+eNE78g8nQbNABc3FlqjvFks1lhcSj5IbcTwD7q9sUuZ7+BmEJpJquCJkY5XC3
A0TV31zWtSilPWPt6iRJJHwJzOHXY9APGDp6D4oKcwQBJSWMbD4dKLq/bYDET7Bb
CO4LEg0SZJmpvSu8xMl84EgL/P6BlU/3XEm9WZyVjTtVM5uvQsK4nscydZmly6Fc
Zt8yBLMN4+ozVB8Wj8lFiu96HNMa1pnL245irTvACQnsDQJMPjScMilll/DZ5JBC
1hZb08AqIhFXdgoUKW/bXWJvNRl+GPP+d/ArCkO/XUKfYb+N8kdebLc1iKNekQQD
4X/IIfKBPSSZoLhaRBOD6a0KAh9ocIG6BGBeBTOTU4P/9EL5lSNxrREjUwn/R7/g
gKyIsk7K5orNhvDcJdp8R6sj1hOolXR7QA2pBRJ9g5crFHkjjC4Mn1sZUEqPLF+l
xJDaVI2z4NlUnyaDrzyYzHOhCTtHTvtAFDPAvlJZnBoRjt+p/guFU4RRG0gPVU6Q
nsWpfR2mnpTHn2jSbFXMh83SmeiqG1pghVgeFdH6vG6HUYkP16+Fi1NhxgNlTE/X
LoNpKQNE5t/KcFsetn0Yv26MGM0jmersHVncCdBmbSziNsSi/YoCEyfDayWYpkUB
rcJIF5c2KCKo/Moph0ocNALPFtohR+nwHd04n0zVnpBxtcFB+JjOaQkDj2g80gLT
Z0BFmfhE33vkrqSpVIt7XIRrEtmiSbEpWLxCLPvjcUoRhf6zn9m6LN9HSRZdbhJS
LzkcFSgrtQU6w+AT6sCwE4r8wJVbyziKpW8b7ta+07b2KaIdG+aYXCIi0la61jqM
Gi9xfAS0GgffKrXeoDQqqRK2Djr5NZSUBfOp+GWG3oxVCxaSKPn5yrFVE16Mpw0L
kFx0UQZnXV1Mc23wuDT7GOLf+HQmnI6OhhZSae8YolIhWCthETE5K1iy5qd+Yx4/
KAu29t2rCbqN9g6B8owRFoFD3VnoTwUGbRp+sSVQwdmXpkI5J/c5FDyYnP/IUtOX
i8IKWNq/J3n2grIlddehn4tl/fD/Wpi09nO2Ai/wTOy0aOhRQ7R52JCAF2KHTGBi
qGN98Frge9N3y3Kl6mnkc5GKkjVgNN1BSJTHFvR4MqXWgewsK7+sGZrvx3tShY6y
nr188qE7idqbBC3zHJYqn2SC28kK0eH+l6MSgVJO1GhJ1R7BM/MtNjujCNaK3g7z
fdzFEIB1154gU1nNuc9jSS25EO5AF2MWSey+4dEq1Qi+TdjIw+TBIuRDI565th3W
AgVCKyVK5DiqrOAfwY/+eTd0Y4oJrDWEhv/Qe0RbavRcrD1zjytVMkuFo3/M5kk5
QqbiM5adFqv518MBX1YoCOoj29q41NopXcH8eu8Bi7BsCTf3pW8h4KbowcSkP2WU
ahk4f4JoAW1TuKVJHgDz0KKynzd15W5PJxKldIOn0/LogVutK8JA/EMlpSHju+Il
EUSqoVcytzbDd3vmaAlxMIb0266c2rPHZsLV5I67uQT3EMTicozJsucqHkysxny9
Om0SUnRsWZ8xblkdIZa/I4+qOYfgK5M3Qw1ERU4CPmJb/rrJfkjIP46mrobHBYum
qcElyAbMFPz4HDDZ1c7WfX6a9wLR6Rx/bMMEvicagqac8IVap5H23v7ZuNeuq5Ut
VAtvzkFGZIXusRy44RCpPis8XG0YgPNXVLChXNQaqOzE9hz8NCHjlxuXZElxNliZ
Twk10n2VmE/RtrwGtShhoUjEILEoY1hP4/lsZT5wnQZm60ng0svjUioOV3qH0w2u
ALaspNOB5HekBn9w5osf1DrYhy7Mw0A9yuy2Ors25DoaZfzgP4mL05+veh3AAqXg
9Vv/iH4BC1g6XAetExolDj4VzqfdrGTljeyk5oy+pcKOozZXSZBCG61gHWWGi2LN
M1l5nFqanMwa3EHdIApa4JjE9l46YsbWfCl+p6SkEaaqGQaSgC2ipY8yBfOsjWgD
DZ0ocurmL2a6vJdxzQxp1DVcWYZ6bIhsrySJm0XViPpyuWOqC6Iqq5i/Z1lLndBY
4AfOm7yFfPCBM7BTEWZrIJa573JBe/8V0tM3nj3dSK7d0gJK0GxL4fMMEBipCqnJ
xi4svWhxxbhQ1MfduuXV1swzDXVaYdTVKCPHafMU7FOL7a+AF1s5VmjODAww3kRc
2OvtdChvAzX09zby8+hrX9XvIjxyLCaBgN+0Cfzs8Qcj/66EC4Kx2aeLxZYg5zZ6
JVUQTat3Jz/uHnHPwRPLC/40Ag+9/7iGK/4mn+hdWEk7tt9CsBDMY8Ok68S3JvdM
PDs9ztobtmFjwZC/3mClwuJNBhuRLHiWh5NskRRekzn2j4aQj4ChSUdpYDUbUAGO
/5wdPRl84HvlxiP7B7tCwDPGL6hxy2f8Nugu02u9XQ6Dt9CbxiVakt84b0wFktr2
6fgjSAjRkkSWBljghqx5Rm3I3PbL84XADoVGCwk0bfFwzsJhaOrTk85JbXQuXqxC
4e6ChIz4leUkNzUSfYxvlaTpRjkXqDNLlUti3CzfigTAtMU6VJH+0ZxaNz8D0cRk
AVryzIxBYwhA8BV4d9Aa0Scf3jHuFr2MnCZ/UiXQ+cwqHEexSSP4yoIWY5onZ8hc
U5BSNKhpRwvVxyX9rde05HDuP7vyOh1boyjBXRFrrHj8DOEs8us18ET7dnZ+zKkc
EtLUcj3yuHeKk1txBwILkmkecJFRX0m6VsHEBWeQF+Lr+EyF2yqa9XL3KrmXKhng
bY6dAmAqEcCUvbNHoryLC7x98NiY0jy0pUbtCVU3Gifi62224PIS2/CAPQusZROi
bwf4tDUCOl1hkRTkNn0rfpngOz9/nz2sUWM+ejRPD+TQ6G/KbcSojEnp5DMovaZm
125OgO0vOnrBy2Bvpt5Plm5x3t/qp+IAhHONJEDhSUmTZKYlzdMB+5c0PGTyNYos
WpTec+FphzU2en2+52C5//dR9F6M/nuXvW0TWjw1PGgCzkTl38GucJ4hbh6+E+CO
KmmzSZOIZ4MU+1otK1iFLkAb2X0BPAsgheS12nYlakVH+wTVEPovl4ifJARbvssF
uYj+DDWqKs9TN+TV/+QFKYFBaXVRxxjyLRdkPpsLuwcxLm4r1cbbnItCRblGuwZo
/7U/z4LAerxiw5+HekOc5uQgTZ+jVj3SKvmc52nOUnZjp+EpnzOE0ebqI+AeLxxh
LRC1Hl6nzMjlqnhGLrBBjSRPDVpFe4ErSTWbJRqUB/chwTm4kcLDU0lN2u8W3ELz
F7GESOF8ICCHFH+4Z8IFw0mXgT34Jx6r/LOdN9Wv8hUujB9C/l7X2KqEYb36d+Sy
FQ3n4Su0jV8HgEgsWYyBqPpX8iXT2pM1DMir6MgDwNm2Y/WrLgGkoWYjBrT1pw19
izsr3jPgE0fNPoO5ywc5iXGA3J54Z/iydC88M3RL+QIw6Ei9smUTMUtGBQ5D9Pwl
QNeX7jVl0vFyKDw827hNG2g2BDwJwhP0Sprz+yh8Qvdqv59yFi89SZbjrPpzdR/A
pa2S45XSZNGNLWZNnm9mhaDzi0a7TAmgB2UEBuK0RsOf+XGCeHYTTgk5FyHVZiMR
Hasuj9jWi6ReL3nVtjXlLBRtYz1DJd74wrB1euffE8ZKm11Gg4bU9bgsPCOWRfvN
GpYqP7EdG4roDL8N8aGRno349Xsb+3JBSMNDrR4M3dJVOF3V2+VU4s6E+tQnDW4u
kuPsfy2whA/eXbEWMgAzoW8jfTgXDK0styd5gKXznc7pzSA0vlDLupAFmJ/Xm8eV
UeQ44gf9pJmR123R3sI/mxHqx3lMhcH9+xZg4Mjwm0amQGLeh3rJUFTZ/+n9HKPX
vs+JMkwuceejqMEd+vQKWmgO1SK6n6pfpaggI0a9uuWefyzrFi5L7qIQA1yQKjXW
YwTC1GtAnhSZ+dka48C6wlUXMF6j9rh5WLA7381hfwfdYDd/qfjg9pB2hWBbfNQM
Ruw9zUggpndsDF7QmBTUD3Ba3xUNdtDRhZMCQ++JUdItgNGYM9R7TvcYX36K0lER
2vXMhemLxcP4y6hO8EC2oO9+/UIRmSYKyMTfBP0rov7FSKQo7ka3g8pLi3zdfNht
AztfK+ZgZEUz7PEdL5aIC78llTDXXQ772ODoqzlWX67YFu3Nfj7/GMyMfKWDQBeO
dIEyP4MaRwtFOPiD28Zhkl3BznbPBJfoWTMUL0fuF2jciP4ZrsL+AxW8HMGjfLmX
NtAP6emNWD1jbhtDU3SaQfQxYHB/XYFOlm4PeRbkvEECoPg3GWycVEL0A3JeKHbU
cKWHY7h7QTE3D7XDa7PUSi2ih6SZ5nrYCAhz3BjYfnKe4tHTuoM/DQF7p7pbmVZX
zK7cud0VjSo8m9FflIPJlOFCQtuZreUb5f9WZjrpsOlO4/KQYArsCZdSEcjc1wiS
fX4upNDjoTx67rPsP6HWElNCXvUuVm1Ks6vFU7THI4PT7h1bnTWMW25clypbUmH4
kLtFqefXpp2m61TbrQWepiUVfAOmxV/j+izFqTjB2G5hUc4WG3jkV9ViRSmIksYF
uYap33+6IKZ5mAidaaIKTm5etFMqbKTEekzrt26hO49BX2SVU/aUkfWZ3/zBOX3W
lOmSgnkEBdsPD6wx4Ml0CKBVhg7FyqnB1lxNC6dyuqGEcpItr2QFjKIKg/P4Bq6T
00CIaicv7SMyKLxFsu8LJpnXwV2xCXk94difxIpeD5Oj05BIZhb15BqZwUYs+ZK+
IwYr7GmviswTzB2sTttF0ujE7yHnoTpY/hNh1idKveLe5UXfF2+E2qqPu/bqsrSM
l/ye1DQOVPOu1IbUxQp8xkuCRnl6GkfsvPKpnwkHWa2C/LAeA9B1cmr0nJcXMrWM
kWPAkrZebXXKlmJWWObjAOeu6YvE/hbGlTBoB4tsEhgrFfYGUk5ZqADZAES7k8p2
pxnE7enkFWu0Baml8uuwiQLZC7rtgnmGd7k3WhONTHv3uD1ucVedCes/g0DIeWiT
yRf0qQe3Jewe3H8R7fAHIZYsywX9Z6PchrVhlItJLKinWWtJ/GhAWI9c5qFn6Wzy
+iUxVRhMRtn3W1ROZq86FTygVKaq8T59JE1DqcSls9kKJGdwTn1XX4DgLr6HMK/6
8+cM4fkoELO8/CzQx635rcW5JbwM7D0bKfBWpK9zL3HdR3U3vFlRBzArL+lW6i8y
/jpzJOnZVZumw67OUXPi44SdzIfohiKicWu9jrh8InPVV1bir6snMDBKdPKD/vRE
bMIwQuaFn2RW0N+OUI/hJ3W9I4tuVHhIM4Rg1bSmH2x+QKzAMtpLClDtX61ttS2L
xJ/iLgD5xxnlWgM+14BpXipFFEMmuXHpRQm/vb4UqQs9SetfcjWqPv8sU6sVGkyv
PGczUsE+1lhamrmW051c8wq3XgCR7r7XMgnaNZtzEdMXLlrynzTSEd6fNPDP6r97
672tm1LcffBnn6qtjSKlWe68HDxBxLUJmznZ21QZAf72lBMR1EBvtcaUjXfKMUan
5YQTr9fl0BsklVy28wo26eZdvwTIDDgP3YPdAJHjNu8zkXpjye4ASSsI+eClmMrA
wCosxHePbIA93uUQmWAbgkUZJCzJ8StNkXGlRQoBUIX24gRVD52aYHLPQQfpwep9
WN6jm1h96pWNaKlO3Xt8e7S5WAmuk7yNKgmnkeLDjuXQMVm5hn6Uj7wj8hsoflQO
Ah2fHQxuKma3CDF0b+GzR5DeWOIUOZj2ha733b0X82wOWOzi9DYe1YqiDWIJF8Qu
5LD7cZo//DFvU66oYQqpQg9cEHxXDUFbQbs3PzBbnkrf7N/E5lWM7BJVQmIlTuTy
LfR6w3c9YyGB21CDNikOhdQ2CJ4jRPUB48KNIk7+KkqA2s8lxHMrF9jYaVSV/uwR
cE37V7Exk34C1rpLxuryvUN2rz4bVTnkwm6mPbHB9q7/Za9lcNLqMJSYvIHwq0oz
SeC1rXNGtNk+Of1W+kYgZ1v0FfE8WeSOfl5hyxjG5NzGZBDh0uXoVXIZ9D7Jn5Cq
ZC2hOJ87tITQKeBjt33AHp0OvAUVAIMSW5xjqE4uRzhLXdNk38PPiRB+fLBi0W9L
TZw8UZJtqU3FHIjM6QgQO+LniuiXg64oobYjk+DZ6+GCc7dwr3rTUgCSmPZBNND9
rOaOLwBRg77la53kx7g+ok8LEdzG2JDJyVC7DymptgzaPO8Lcjd2Y0hspnzFOJN8
+h3er16oxkFoZIanJJqkVCBSe4ovhevuTWaokzSQPpD8L0KVc3zhF4Kwb/DIsTf4
ZigjatSwuuZvHXZQzVPNZ01e4YY9LFmwbArP932XWkcT6Irds4J0qtUSdsFBbkK7
XY0SWzDD+UvQMPuALSDxeyGXkVLHEtgKvcQil3I4GLCoixYHf9tVzQ0QRROrtNbb
xQ/phZ/mekyhP9qAHUNrtvl70U7Q6N9fLi48vp8has0XV7fLFcCg6IVseGMIr+Vi
KJZsFw/igaLeMFYVTG60/2XoUimIzhNfeQsH53+Et7BXw/A5Pi7Ifc3Vdy/WCk3l
5Pd2BhWn1FcEQ6xO/xfZvu1+DWNEbfWkhc6Rg8gFk7wadvaRGN2FScqoJ1amEFrh
P2TLS6lSQ9geQO4QanFUqhQ5f/K6LixAH3F69GDWdp1OjjYApcCCKiYySugexipm
v/CjacptBeicRylIGDhASoEAzTTjoGwF+1rXr/Y3wxggTTNq+CmjLrOvGkxs0C/o
g5MqIAW0qVUyN5KGNmyB3Id8jtc/Lcp5HpicRIB3zsTxfMxfWfpztFLsAPdWaxs6
ue2Flz9K3z0WkIlfUZpIhBTXgNtfCK8PbhMNmmJAqpfxRq9Hx6wm94GnDMSYwNQz
UqT7e9HRxs1ueBrxcJhW763zBaHbF9NeY/lMFO0TEqLGb36OWeYRoCnaDNQEfr0b
wkYeZpvtYqdtqybWwTrnC4uGrphSq9ym5g3HNVTCAf2Z9QoREzQhnE0IBuukbm1A
8DRHx4+urd3cFIP++8b7B5txyQtPFyOIH7lYDqAoUCDQqwWXs6E1TGlKd0V1XI2w
HPP527QJdWfx7a1x62scqsBkU4L1it3mbEUj218QN+tuNTaVURu8f7cCEk3QRqsc
RFbh+iGafma/nHy8jyxXyzF1b2UIGWIsnFH4fI21dZlxc7sWCQwFIjLOyfSDRVKx
Yq7re/e1oqbivOo8iLzFeiB/p4fTrwxjb136VlhwSdRVRGp79niUgFoQQaeZMl17
j8zgk6xGzJR0G9O1eN63BhCEpovKVfKaKL7637HjJjx1PAsCKfVuNmk3loavYrXV
tZyktpdE7bg9AVlrvzzTwvN1Nq0i0QQSRZ0EKqH9NkfW6UIvuj2IS7NH/TCZZhy9
KGYa/R/a220mdXSaiCZXRRYIlUiXFyHQezU5DwQmqXkMnrRq43pU8mG2j5L9h8XW
9yE8UYSne4y3DSxUYmPoftIh4EOJt/eRBRpUyr2RDw95J2kWnodz6kamXw37uQQu
effFXVL43FXJrVmA6AvbjnYB4Bm/I9psWeMg7YIbDrynqdGFK5zvseuC7NrD9A+7
0DS0amZ3jwOeYKs0V/x4PsUt/b7OTvSXN5ngelw2sCEfICGuX0NLYcBOCIvW4A6+
7YJXekAge+Qi67p+lU4umH/p8T5QxgKnRkkhzRsQVMMe06eK3/HErYb33yDtTBDo
7szwwEdp/9uf4dKUy5tVLa2qsxQRRUIuDoQBBn6vvkUmh82xPC7aYzl+wOAErzpa
uR+dK/rXfLPj1n74NJf6mKm44VvY6cUFdqxqfLu1pak1X4xpuDz/8t/+/80FvtKZ
YogCaioPdq1eL2YddMTA9+Rdzw/8vtf0gR5sSFUh2UXh2V+lSzlbqjr02rnPxzdf
KUNIOHnlcQCDxINRy93+LIkLmsiFoMJ6FXplJKLN9GvulmRW/wU+4xJU0iC0681B
xWHySsYTYL86F9/QQut2m8VgV9JezR3FmQiT0my3S86IA0XTCJ11miOMU/7LNE9y
/mGkpyitPf1xuOvcwph5dyuAJYAd+rWvmStnv1KAlXE+jN1WGL25E67yZYsDreTZ
BVpsu1vFD1zZbeVwIdi8fZYWwx3XkAAsgJ3FIyt4EDVZfj5cn3Z+3xHsrr1jumLm
bqO0V9sXLLGrkjI4N/Hx3nMlmRWxjagFCSlKiXYx07GVepn16ymlsLIPyFV41pxX
CtUv7K8eMVDdN49JSLIvJYvBXBwxpkBrTYGFs1DTd5Kt4YmBOnv9jHjzMPdGBp1N
siPQxLjfidexfZYOOWFQ9aO2RBN9XRP4oWHum4MZvr4W2IVnJQmrhbDT275OFutg
B5KGewdC4iGFfMlUMQM6Pl0kFYJTSuXuEaqueaq0bHTt6huWW7quKB15qvatkNyU
8DneSjOQDO0JwJXp2GUbRm5u2m2hECl+Qii/cQlHWw5WBmBtE4Mh0ufcpu4dNl61
eoIpy9UnJPI6BEQemTmGKFMHULcsD84vsiBXAme0u5zFY7yVLl0/Sfg1dhnoHMVV
B5OhHLEcDrobYs2GW/uNVDK9c19gZzjOUBefEJfFuuzi/3p/ujiICYMcIGjUHTjz
HBLlpz3mQ9vYQzFe1zor0/1PcjHWokXOIqO/6koAZ9lx2scUd6dqLnzrh6Y4HnWh
Qbad3jbBo8VT5f0bZymEo9CGWx6wreKTUj5dTV+y7S2OpMDf0uI70Sucu/70I0m8
/K+Vy/vKNwzqZSygHAWqXIoUKHLNzBOMtxd/uc2qjhiyjDtO8tnWEUtXeL+63wUX
/yo2CeikVWhV4k5txIf1VfE2zAZT0DwyG4/joqaTsNuRKZfncf4uVZY930a8NVwM
VPm47L0jXoKgNIaJ9hqsOWAwqpTFzY+N2j7uN2hx9OZBkrLjkoX7d1R7Apaodn1l
PCTo7p89ZmMTSPnXM+0WzLbVkWzQKOlsXGMJzi23qnR+l5IaPF/uYje/liSl1ER/
9i48lemJw/IMuvAiZh9ufMSpM4U9MsM7hW5lHPsPoEqsQZTRw9eixQrQpI7p1hc6
3GySFRSrx9qNqPKTHioqE8f+VyHkKwqQpvd7ARPmovnYp/H2qsu/KA7r+BcMv7+d
smsqz7BkozHqdD64ZS8wF56yO5qYaAgmW1Q49ZEOq9ENgLVoCYnkrAQPBoimtzRl
t3Y5AEbBQoilU1OsXwazkboVMsIKjkxH321Pqp+4+LkjTZVPPiPItUyu/T0BzkVj
ZU9IUzRmy9nSI9xOjmod20tGrhJAIkE5fYk7hBnVpQZEgtIJlRwO2rWnrjIlJkdy
bViEnfeMLmJ4RA34FHO6gtXlgk+EjCAKiHv1+4qmHg3yW3AfiErg7qiP5S26TUrD
yw278bTf4EZ+2o/nQTd6N163JWtGCKAL8YK95tqaBb0J5hDzmLtzBTx+XBb7urmk
GvaWhhs9eN/k36ii/7YFILESef+psu8YHbbff0ibIl0aHndjbz4Ns6P6CNgY7UN8
ZuMRQSS38+M+sfAKzU6wr/qbCaMF/7DUCohLtQ3jAh5l1MqBj+/bI+oXiQ7RUUob
pjRqqlQ7Xbs4woTaPILUiMZPEigyQvwPunTrwdIwocoIwnR6DVzJliI8ODB+WFO7
4ORkPUf5Q/Zc4ykrsnavw/TLhW4tN0wRojqb5zQHUdmQsjeBdc4Tuu75PD69pCMs
Je8xmKngc3CktTyQVIzQmdYvzdt3liXIzkSLwc1poLeauw0HerFoi/g7NltTxF20
H8DYZHNLu/9c1/07x74ADqJO1fxQZBJJ8qSKMT19KPBiKf0E/+aSOMKfJR4isrRy
OUdt74Ovu0qGUIqoIU0cHf1XsH/aWqn7jdoDqNMq3QmC4CxDVa6QsDasFkfIbplH
2sTeoZbgg9tc/sfYv1U2YNtV2VWwaQqeW0Kzy2Tr1VI9EULajXKiEVZ4LFRtwccg
y2v8nAjoICU+2V2RhSRdryeHXk39o1m0quIRIVaILHsXlZ1YFeOW0ATpaAF7c7Qq
YwXOBky9fa6gMVex+N7nCEqAU82fnGSNas5mnUrmL4gqZ/SGM28cCnTzbdeTl1yl
H2eSYOpC+Z8zFlJ7+EsqbfIs1CxGCGTVlrmc16Xoqf5J58ZEn3p3qVVVua3PeCE1
GlH4gkADnKcZqZ83pC+X8POSrGllbXAHMnXM2CCLZvup9+FCHEzJPmeF/rAza9ye
raFywaNKdQ8IK9SfJXQ4mxogjvjc0gX9GTKJESnvZKxxc2z8XL7a5iRyBwYejWkk
LjEKRP1PoE1EhqGPWavDTZp/Q7Ug2p8CoJPisV+/NIfCnVrI0qx0kvyPEzVRB3tA
RuOzbSgexm5Yta33PIsEDBmTBY9lYaYicmFrwKvSJQi7qV16qlQRe//A7cCBiOnc
PAom05rjyaydj6H/a4hvrBGX19fByMKe0X6jBJNx9KXrL8lV1J5afs2IgEuAxQPr
7NSmbS4IeRz990BgjhK1txqr9whF+oP2TfJF1BdSLfrPIg+EM5eInrdAS1Q8Fblc
h3XT85ogH48ki7OVGqlkgMwS9K3LvwIFUR+DL1LeB1PUfBfFwOBXjeSwtfhkaT19
lwVwPnkVK8UB5Iy55tu6mwkrXlguy1wmPI3BMiZlOmSxxr0gaKEV3TuI6bTk7bro
rWYwl5yOVQpY4So7yuumas4q3PHVKy7wHUshRv2HsVoQCPsR5/TO4Pv6R0Jfe/J9
VsR3opuusLiOno60H+AmKOndM2gVUYfuqAp9yHsyaO4Zxhylu7pXt9LF93tudKB6
0qnj/W3rPluZIGkVZCapQnaQrhfMG5hbqFTie0KkibMmGARvtGEqJr6jbiYCZF5k
v3VV/V+0RAXYc1c380YSHXHOMxPiV4JCQziAkHMpf6X+kZD6jBt76Z3noYpqCnNr
r3rDy3mJsMDNrv9mwGjtUgEjFbPQG166OiI5+aYViRNRo/oNIl4FY5J4uNyPZtS1
mjNxwzRc/3cBmYXB8s49rg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JCA55lcKphIwV6T4yFaahbpvxxxKyeylAsRmPzbbGNlfdX0HBymABvOiIzEAS10F
wQs91Nqdwfg3GUi/4Mkiw2JY1uo7dDSx+9EXmVQVFZNJz/zJ7nePv1uScKmaVr8X
AhT/t9Ap2QkWY3lYE6Gel+jYCykV/BMxXU+2oyrw894lZoYDdU19uFn4ypDvpe/d
m8lcESiyuxdEbm5/QRqGU5PriWt8XEr2lhYy9YhMGRJKekFbFrhhQHf2VYTGyD4T
HhzxT7mrlw606nIvlG0WDdWhhA/y8n+WYsR3ivdQBo3UGi5MR2CmxkbIPv+/cEU+
fFYUCW6fbeoLE5URzvCOoQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 27168 )
`pragma protect data_block
ZDuz0bZ0pekPzJv2YEwI7pRYgMiXHGR5mrnwOW6aIZjLaJzxdO+RBHeGMJQP+3uK
DOqz7kuQdnmd4ezKrvjhVumS29NCQrRlveNCv/1R9E17KqLaK3hxTw51RlkvgSg+
OvE79Pxy2rnYZ3lEOtV92o6VdZ02qhiS4qyivXcMhY2KjxQRI+4TW/3yf69HFeOq
GtsawlUPjlUGwDJmaqmCJbjdrSgTDwo3EczDWLOt3pkQG2IqNSLtZl+r9zuN9MBN
DSIZZEtE3Bj60HZ34ocCqjhGXW/AtURHV/2GBt4eSOkO6lKsOCD1SDH2iwAUoQCD
ePeNkVR8Dp3Yv0wdPX5gK1/9DgWkIhFMkv1gJA5eP9qC4Ylny8CNuJBrG2Xat5Jy
ONk7SuNePi+/VA2jAXnTNy6vSDI1Wn6KHxkM9uCKb/tZ7wJBNHIBf4ieopeNJjcx
ZXVcURjBBiawauahd1fbu4YEeXF17+sUvDFplS3MhS7D9iQSh/PyqrEq6YtBkFYl
1eObb+SAJyIBDtTo/Fju911BoKDZKIcfXu0L0O67w5ewegtcEo90OKM8vf0R5TEq
19ityrQFPf5qvx8K8RMkpnYCdCICBtWHQ/wDyMIOzFUIp/Nuxbfd+dN4wglBf7wd
gjpwQT95nw7IdFR2Q+46q2lCltTj2AhHKh16T2ZBX/89QYJSXNn+uJTRJOq92nkJ
5DJcMgwP8QhQn+1xc6Ly6/MVlTqsOq5ohLeWxahmPSLljYX5tU1FcJb0da5rB/qU
IddE0T6D7RuzXszvtELmwdDOyKuDjbqw1odvh1XNSkDf0bAHSsupUp0B6LbTVYw8
CEeleAx2O1FPe2vRXyp5AqW8lC85c3WjE6fy0i+QLdmqxaKMdFahjSCpOSq5c2Mz
eLX6GlgK6GRaUBbL2e/AqXO1xPkHSZYyLMkAqbDYXfkvzoNvrz22uaJslq4+tzcg
fddZYf0oNPpTdrWsNIGifOQ12zdtfPksft23kozUXEWBpBe0ckxeGydSqIKhsY/u
qYBBV2vk9MvYI5d5AZH2zaSFbqFbZLA9MdbqD06wV/C6OY78oHN7TuifhXhPK2Km
exazbZEHwpI6owa25wGLpY+131XRfUwvw7DG6O8HcVFQn+h9w/JXQcL6TsSFhryJ
Tv+VYRyZEGXAhZjN3rytkiGVyDHxM5n0zUieib1iWaV6gTz9TftH3IetfqRpeEWc
TW2P00gEj+MnmZ1Y2Ri7ywXqP+SmJrLK5dwGKp0qIOvvYVLOPSxrFlLkobsvunsL
VVlgD2raDmE7lHiSJfZ7C7y4kUvj2Bx+0+2i/c1wjbZSWw+ZAArDfQ1EqfOqA/5y
TL5ZeKZAAekrgIOm2H1Jcz4OjXHUrHf8/rMZuO8+xKTuOQp9IUWFxOuEdwqjiDBv
2lI59C03fTLXOGtyc86P0fzaSFU+qMml0ix2dZjh3mhLAC3hmNpOsNSgMW+CGr0s
rbYEjhviYuMG73Oup8hC4auRrafAtK1ZSHdE6+b/oIhbSHikGsWIJNhdHt4FyYdV
kFtwoihMw7XP04VAlabdAn2WyvO5ZgHURkpJzx66JzQTfs9bArBRGW2nMmkKHCDo
MOiCcVaCi4qHuw5Dl0yp5eHIQVREsIOfzAQ0o6f3rLA7kCWft+4vKsp60vy+93pD
e/0UNxVAYnxAmdRRpCzs1CxRoFwilFxdFcO4ziFYt1vQ12IxoBtw5znY9uuZG0cP
Tpsk4rkh+8LZISPs4h4sEt85Zsgmh6xM3sU4+57xTCMWnzc2Z2gy1edgwn1Yi0ej
w6NNYqV+wcJp65DDdPr5AJ/+LTSkhoFZVtMXOGHwx5Y0sIRLAJzYLrxB0i8RZUZ4
vfjGxsMFHagn/MfCCYvjsFP4qCwdHpumZqle+98Fo6TZIyXqe7fdokP5RBCEtzvC
q412Uuo0UdtO5ClsStgsZ2ydhOPQXQb7+uritqqHUFAugIcVMF0NT/Gt/iRPnWU3
mycZ4O6RZ0Pd+L5teOixmwTWrSzEcuSRUUXcBFd7ctAsMtio/1QKoh0xnGJNjUAa
btQ8KowCtZyWkttjJFn+2vTEd5qosA/2vc8vNl2Ya0xjXS7XIpVAx3BhN5VJh2gz
XjMEQpxRH+B3c3TVV5IC1Bnw6Vj4vY2igI84Ms8yIwdG341R0ER5b0EKdSY00Dxm
MV320QQQwOZfXQ70lLOHRN3OSwP5lQ7j2oG/9O+kiKvSRp5BO0KMhW3eQfJwZFbW
vDd504UiUr/qktPOdpyQBM2XYf472OKHXycGNMZgBMfvmPWwFW0vWKyjT2zWzZlv
+KkmEOTDuKan4qfXSeAU6nRIF2plxNv6zFyfb8TqC1cauy6Vi5l7ByE1wGf9tdjq
qxN9JE7DXwSytZJqUnJMjnN7wERTLpiaS2oxf6rU8mDzmr9/FUlA9Q2CaP060pML
mKlH2gjzPSTxzcS2149Kpql/SJ/WRW9XH4Pj9/Ne6VOaaTC/cITTLt6qyT88ElfQ
T3xhFSWsJallc+KWOtYmVM2XZ4VSEG56R2aoq4Jl1y9qLXFKOtBeGf7Tx0bGe+iQ
rF+0U2el0hEarU0n+os/+pBD0HdiljvKcMFH570tH5iFO+exCRwB18xsuiBqef/C
0tmVqSR9rmxMXMLzy1Ef1HrEq5yNRhnR61Zd3oYdxBAt8Ix2nKS9LvG8cWKh7NHq
b602IHiQw/Xza/2kZF1KIenirdr/0mzBnmTxynJ+YiQideNh9rjoCNXAnGY52StF
GqMLLfP0N6xxI4FcdzbbieXNQj35lnrLjReDtaLcgpj4t/E1MR8EfL7q8mHpA/eQ
Oyul2HqEOx2XN+G6CMlyk1hJu1+0cM+TKdC/kGLEF2TGhk7mJbI0ddg0h3UhOeuK
SbehtwwKxryOddNSG6w1/IrtN0mgysPPqs2ZbB+4P1pe2p21osmnIxBPbQL6DA+5
ettzIj3sKv2bqSz+6pwGzEUw0eUS/+UJa7CPts4Xfxwmj1TxkGSNDR9sYm+yiYAA
x7Zs4511pgnZVNolxu6fCFIrdRHa9zkBHxFlw9dthu5KEpWli/CWCkxdmyl5ki2/
f297j3UP0gcTeURlSo1XhdrjFt3mHt/OqClLaFKV7WIgAWJ6QSCPHLzHDfAS2OdR
fl/dUUxIcuIcXHM7GlQHNSFI7uXjekiLtHZo7RHj3zAnxDwH9OwjhAfd4NtqkQCZ
GxoXzCPza61tOdb35A0E+nbF+3pAj5jsOBhp2Ern29+jMF7LR0gl3XZO3EqBAdrC
MyaixyhOANmSAd1csLWDijmbKhG+GmzYS53kJTUkfA+4lfvN+lYdYpqMIG7o/zMn
Djm9qRoDSLJz7u44/2J5+mojmExSULfwU6bSUg2KCPBQavDT9XltRdU1qoaK3rMZ
Pjh6yytDgTaNYVVVR+khRjilz1yr4X9D66nLfV98eVrpHThHK/wDY6uEPrW2fKTd
ZSwzdY9FbBH39MovdKPueZDq7WTAGgGJPB1gxECFCbJcUZXXtpZ2gT/YG0reGW1s
d38cznW63rkTgIwtKrnHswyNKz/J5qpkgcZNyjN7SFSBVvcEeLXQCSptZYSLVnGz
GEB6l0tTauEU96X3zIojUD/PvV/tMDOTpfvZrCPqhrxUceZkMKbdEYk4gQOqSmVV
gYoxH7Hvrduc9kn5Zf9EWK3epwOVJXWF7wN9oju9ya/oX78lbZOO/leFNDTsduTU
2cvJUmcCY+9Af5fBvsPOpg1KV0s6y8QpatdK8vKA8U8DylxxvaKGmq6aCFD6+F7k
Z+PcJdiqDafD5ilO/WbQ/PCOdOb4qSRDdbv0XBN+lM9V5xdUC+k8WRfwBOzN4Ko7
ijk20KYCEzU+taXXtny8OdwtU3qSIGROLOLbqKNRor4YmF3Ng8xJ5BPemfxLwxic
s4v/9po61csVA9Q9qz2LCUPVkEm1IhOWQNf9ILXJunti8LT9fDxfenc5qva5Lkuk
eJMXIjX3kVJFTA2UTt8dr0z69yW5B0kJjs/+SuVyzxHZaQszvF1hx1b1RIdnXrP5
0Qt9F29+0LcnrTs+ISd08fi9A6B/kss26heasab6x8ByswgTjF2gXmnTb1tAbKzD
F7bGBMOEAqCmvhVjoxFqxQtOf+JkEBi67vnwVHX0L/kwFAu+CPmA5xw5Ykm+wrN2
6uxfaxKZKe9SHWGxW+81KbRqVLmtNp6hXk0/0MS8TdDLFUFrwRqq528gMvuBNQ1s
+q3oTAybAboPdRfYV91YzlYrxicTzYmYVwj/FthoUf8hDvoGz6ecTRVZ1pR1D2Ew
HSxpL+bj98SD7dHurxlhTZA2G8AulLZwfIuAg02yN3Q4raAZ504XLO5161FLZdsL
P0sQ+VCCnVo0bK8riUxq036X1pEXpM4u72K5yE4iJLf4fiPuBRtFLW9iLJdgQ8DR
HxP9vVtCMJ52MkSEjPbu6wid1uRRs0uAia7kiU0JyeNSSe8NLAVXKV6x/EN1pkro
N+QjiPwfrI7pBxFlFQxTVJSuQGB2FNnotaNmzfUShbJJ64QuluTz5kznIEhFbg/5
I/y3QkXRxOLqyFkqRdS5Nquu0iRdmM3/PUJE9T6yIJmSysHzJqW5Nb/figfrUr/8
3AC/EwlvlQizf+j5lWOcvYgAg1qOqTQ/FeXliifzIcOeOx9OZZw/V24QT2FulCpu
t76MnIJsczrmCjtnO5zc4aW6lr+CRMMWjZTHNWccjsvdetIlXnOwJHyxgICmQPWZ
ZLvk5GfrgfDmP20EV8/GzUawTByVzE82doty1xzbnNij6MZftFncPKkytGZ4xJ7i
MZpAXfNqA06vhU4yPI8y3cGMTyYARd6AVsM1cUEHgnL5ZmQBfvbxwyfFNUDbS+b4
UVF0aRaIMPy/wSu2tvXjn3+K5GcJu2cOG2l0ZzxmBwXvmp2dbuQ4CPkc33NLqujX
VPPf1B00jnMPJNwHHJr4ASy3fjL0vGknXMd+XjueidVKjtcWmKYP6HXH/vlouXfJ
wcWRxyIyRA7Bc8gaPsua82rW+ijOZWlOGy6kxXZlC1EIAH/XDCrHNMCwo0rBlbFM
VMsQMayalJD0veI6GefQDxUDvObTW7EhnbAy9jylnCBgRESdOTwWYGHmstLtVdbT
2u6UKnO3mHAhAqsPSRwU7oqAjbqfnDIIchKSUxTTU8Izqobsk8enbe9C2aHL3sjw
IfrO6YYUrwtFJDl0CDbGY7ki3PIrLSkfZ77w4HVKyJg1PguUa+2FHR9lJIXty71Y
C/xHsRikw/lbqKVdK58MwbP/KAux6KiPbXcod1P7T0mki0b0QmhftTxIDUvdiLPo
vrbC6tGk3jKFlb02W8CnnkPNh/fNoAE74G28pSGoeOv+AjluDGLryVkDEMbWv/Xj
jU1tnnqVTXYd/V249OcVXzWWf6ZtNSaEmXttjEent7jTD2VqBfYnBm0OV8w87z6j
dYOmeC3wlhPKC0AZbFEwmE0PsjbYnSjTlmhiBRSEJOs7RbMCpX2bCu6jqjXGHmzc
TDxnDtVRnxJyFBzQbMnsFmmUd5HHXs2PPFJ8ADL78SmYu/h9krnaiKLjFpsFabA/
hN5xD6RLCEFX7hQ4GnIt30OWkvIUoR+FZf9g6BdaaQMRv9VofK9ayrKvxNCMOqHO
SUotrfi6PYoTPF0l/pfqwGwU8jA98z4BmGuqiZm5TrtkOWQQ5hAnw2yiz9LN2a88
wKt5cBbzmMGWMQxqqjNga/RQt5ZwPkcIlEmJqho4ERECMkt+h8Lm7RN/PH76ZKkO
SsMfqDlXHMtsk/o079USJExnXJa4o43tjOPosFixBmvgVe4Oh5gwdw/WAfsUwmLH
J16PSZ4KgcwPhTBnHGfULaoNbZRMxKOMdQJVZUNkcTLMbsKXfli+LEWs33EDYhsx
0wyOPlS65czAFJlpX5JOoG5oNfZohlrj4eGeM/19yGoJv8Tt/FXdIr5vqBtfxyUG
375ZhUIuEDnOeVpbXvdJQkeDQOJomo18OOa05DRCr71nt3OClo3WmfqZbqfAjwym
UZEghjQ0b7xiYE6vmE8npHzT0YBLcQDph5Q6Uy0uw/l1snPgM/1hNHFmaa2LFvU3
/xRYYzyJKlD30gG0CaFfph3X8JMy/k4CpK7fjjH0JgYFnLYVlgK/GQODXuNE8wdY
c7zIA0h99yIggRnW7txjisEGCixsNs3LDO8MHhCO+oEm6MIN8bmJuXsFMG3qH2Nq
rv2qCEgwnTWXctPa+6xXT/Jr3VShGecBxvSDMdqSo207H+ItQGNSZumbYbcj/9r5
UJ8Gpmj6XxpgtNc+yumiR2QePBvOqpBOHGIMgB62/NlsXTvfDDc67mO78Z5WDfSb
A/oJJAGMnE2eL3A9FezxkPk8KcBV2OnNgvwZHEw1koya92iuDE9P3oEjGJn9wGBO
JcWF/j/JGUlP7idvtzLutW69SaxrRy9OXlZPt+3l6YmXBZfu1A7DcZ5MRRJaFAQW
bAJfdDNp40IHAbqAUn3pvW1HrS5lZAa6MB8hrgssScM0IQSYtcy0LXfa3h+s2Wl9
7QcqwatANHOPmiyMM7GhmVC/iCYGQUCVDDUO/eDHG1JCHWyLywYQeNJ4KidTSH6M
bj2w98bj0ADkSptzEHuL98BjU8mAsaq92QrpW0bAp7flnDfSSvzYhnUi8Cf8mVDr
auxpBx5Ujm5+LQ3rua8UfuolqhHbMY7s9o3iw8zmsdC8oeGwrwpyj/2tciJV8ofD
el34R2Xxo3iJEs5hrU8fkRCJSbbRa70HMIj4QaVli2mOvksCDyGQHQLFMzANxwch
bBkTpMOSelNUl/BR7LplLFvrRcRBazxfbFaDGWZtky0WOv7eVAmnvQifKuRTvIMt
L/V70LUgRvvsN2tC7nREOoXQQyU09rettnl3zZcUdWPOeFvqDAd/IwlANsyys48G
H/G1jDmmTitaSBPpW1RSAcAEKd8y+HEd/iMV0+0ru1dEtEnJ6AHrkU4sQXB5poeg
+VxsQTibHRIeHTA5hNIOrgv1WhqXgF5I7+b5Fmt6KbohUkwdf6rvrAadlJNlOUPG
1WTerREDq+oSrJjw9QefXSKLRWDIFyRAJ/nnGalJFZYsUEIGG1yppJouJ5drr53t
je44KisXo0Ppx5XlVLmNjld/0rGTYfra6ZhlyDyqxPffy3/BwkaUUUYey82QUM/8
z3Kzgqx8iVisLOiDH0TsYWDM7QIY7GujcwIJjG4s+npOgpVfKUjVkIeT89hreMFq
R1u4ZinaUDHP/alkl2dOXR/8HPnBPFsZ8Rnp+jHO1nfgxLlH9QhuXZ7N2V/rqP3c
gQXjSw0Ut8/kQENLhsDWTCo/uNTBgF1iT8GbbjRovyq68exxTi5eoAq3mKQWgdN4
TuzTyQ4UGR6i1W36DYRzUfvetqTZ/R6zmsyxRq3iSg5SxGxkV/+8N0U8G1H4mB+t
Uhgq6cblkbhikPx/hmT8GlJ5a3Cl8zsHNhXxnuzv5HbumDFbO3Ypsjb0/O/4Ru+m
OQClB2y6IG+uukEdOCkf7j0/lqLaxS8Sio70/+NB/wNpMLXwOfmCus+fiYXoFALY
gds5nXeG6c79AE49ey+cuupJBkIkwj9fvuAQRh3Bxy7hnVnLDnj3hpvk2qf9z4U9
YCxreeR8iA6hTdu+/hkkMG7VowGrlKpTdbTQ2fU3RQAdoiyo5hBJHvnYAmQWK0OO
5YOCchRS00kpOoBVuWbYfChlOC6wSBz5+3T5zD4eD5Mc774wTLL7kumT5CgRXI74
xO4CrgkjuSJcKdBKN6Di+NfQhb5BkJTeGJfD+bJ6LniHlnJbQxTDK2HYkdQTG0Xz
CE4Lw8J85rWtUJopCT6CbOksaKJhECVKJfN/4qxi2mzIf9bQGl/Mu25VELyvqbq8
KyXtrzr67MY4ECMt0eUaBSORlSoNU8ltF0GmUg40RV/U8TzYDAAGbQIAGdgp6q+s
ElEmPX3f9NJFwAYnPe5wW55X5ITaT7dkxn8kGT8dfOqR4KUnJp6hIzSOLLJtv/+z
d3BBLoPPf/lchP0d53T9oVYjIDr/teGcf6IMcfzGVAfvl5EF9wBfbvEN0LGbJfSY
QQkzsKwd/I5CMcIhAcELV+0Vhq2gNX3iT21dUgO5FtwDCTO+yhVOcyyOm1/5LqNS
zlsLWjMNw5k8xO+pfooBQ7YKsD13Jfrm3i1Qb8Ya+k2iAdTH8RYyo4LYnniHCv++
KsBjJbp8O2yxDkFhmWwC+Q2+mz14yPs3yvbbPPJSrmVYLo5Vy5axwt9y44+azm2f
xFNy0Pd/iIsJ2fWfKQSrsH8FCmrYb554AVloX7sC9w/5UUjIId+93weLaRjuhSB5
cDq+yHvEhLM4EYYpjmgLGo79BGzCVExknwJb9BzBMlsmQb3lS7hWhXkKXHGPnh7m
oONW9f74k15IHLqC28awdmyFtP05cc6hT5EAYieNU2mw/SvzVn1wsFnYnTrTclMY
PLwiJDF7VNI0va1cV4UbcwWFB/wjhJXqXIVF2Xcvi7+JHDhywVW4OEy5faiNWLvt
s9upaALSOIeyHJexag6pNglkX+YsVwF/bR0QKteTYAnqPgmqsvAzk0MKoVmPuOzU
Kzm02gwme1dOASyXGmvIpBHVw4y5vF99LNZSs9qivRKUPL3kxP1GDPuL8YafgjOF
o+f5x9zCJ14KkLSoYHSMjKvgw7vqWRtljTGlIL8iD4MgqJWlQrV3n2X/E8PoF+QB
46/HnwIC77cTCdl2L+FecBP5rmuUlv2kH4LCSJvwX7i1rTbmzOffnA6pOxcziWUR
CT9quV5MTPAJvl1zgzY0H3m4yvhfIrzgAABF8i0/ZhOiZQ5nyqSeLOLTImvgInN9
jA3WApEW8OI13buzVv1zTELWwkSA7jJBghuJlut//0f2i0MLPtncTS3aKTOTcuJ7
4hLfCj65VxyifhAfyqTUGbW9LBZUWb+MODLs68qAHehbxUYfo0MAhMyaTOcEE1kK
8XuGThmQ3CzBazUN5ocSr7qUvBwLbD+EbD+/ueD2RWnjeZWBtD14GenKPIkQ7WTC
gfyg054gTDR4I9PJTBrHcUc8At+bxa4gIQeCo79hZn+jDGl3a9TwzTLJ1pqoIbGc
ouSUYS4mGF/i0/bMeisgPHoxSp1DyDoyyjVSiKlv2iV50o4hQcWQl+lSIa7ELKxb
q4rjqXY/NKpmQdlTyFLyw708EqkVcs1uy7nzGjOLYmdT+996/4jtjLJcvgvYyqGn
F6nMIjbkm4LBDMRvFdpiv2g9YhGzoMmxrm0XxzBWNbUN+jiFKQ2ySqw0RkCOit6o
hcWh8A5/NQmC6zlEFoQzMb1YUSs4GEOIDDIWwJggc8/MKTDz+ZpNvozHk9ah/8Rz
yvLxudVxcQG2Ew13Wmn3Hm+aP+ozrz2406rllbPdyXe/yxEaa530w4pHly7QQ1ls
BGJA3GuZ40vL/tEu3xoIEr5GsxhN9ONnJJOnsVCjFvWxzZdOYrKDFFokVNjswI/Q
8SQ3GTN4g6vX2tR7dq7gpxY+poKXT60ByiO1YBySd7BscUrmCGt8fzanKSBD1X5O
RkOHroB5B5KQqlViVGaM1WNn8dADKmMmaVZka2mNGpL0krMw0ZSc0RcZFJVT89Je
pk/pCyIbORqHp+J5u9C6MSEiQxHiuD4rQRUTRBvSbXima9UTLYCSIdhtsXV7F7dL
k6tTdv2oauayZZjYeNqlKAWG7ivmPUWzlJYfMSzMK1kwXJs6mn+bLL44ncVVq+bq
VJarV+Q73h5rUUlo5zpsc0qestIdmBNnXARHrXRX1r4xVRT1oPibGqNzKLN22ft5
E1sQZG4dvkzIk3pYFty4WXu6CtbOm8O2sNRU+ZNtMG/1EnYEi+Wg7R62kZb3JmVs
Sjknk7E7Lm5L3mR4jbtHRDRDUc08cmO50Ah2oiqu35Tl/WXoI1sa5bVFiWM857LX
hS9vHedmTPUQpKm7IykXXXHQ3Ygua91xoWMo1kiDS6aSAYvJNAsXhQxmL5B6/rBI
TBxL0GMeVwdu4g/YrH7JQCWzalR9I4kjJXqlORKUxYEJK+Ag226kWk/hOYwxP0uD
lRiFwJO8jgv2kqmEMi+OBKN4xdCtn0LhSN7ffvsByvPBHrCSj96CiaG56A3PUY/o
iLLUs7tI0YL/a5XcBI17gfq+hUpca18PWBvA5Py1faBT+4Y/R6SZ2bq3M4JKQc86
JQHLEkgH6+pvPCqXLDW+RMC63M+xtiLM026di7ZQGUN44xB67i9WU/WdeVgNpUSK
8CKHObq89smLD6cdOhyoHO2fNe9ufRHAMFZ4g7R7bAfvI639rUFWxn5Yynop1mxy
2EWu/QpCjvhNYtWM5/pcSIk3OIwTlj5d3LGeQvYgcA3Guvj4/Q8L6dMX7TOZR/DZ
jfghp0BJmBvaq2gysH0goVG/9DeTGsgWhDMpYVDnDBklG/PRsFbkLFCfnS1DGy69
0A5xdhOupM2Y5YaJC/iFiO0nErbBjc6JpnR9lo3QTdZr1WlMeizPtSvcLLlOvHHw
VohxQgbU7ebGK7XXVISBniC4Cwf825YzAw1ZoKJ9rj13xiz1ci3L1o92MjlshGkj
s4XY/B0hnDfJOcXwKLUcV+AqnsSZDLQyXt6rU4Ony+Y//AFV8b+/rEogmlOBfr4d
5aoBwxBquH/OBBXDSz7AyWNA0TcW3gDhUY6y3N91TUORHbSg2WkGgwNggFZ2Q//h
hX1WZZvaGupVvxkPPHuBFzD6qccw6Imo8FkGOUdLyGXESe4ul7GRHPjT8sOJwl2q
jaSnyBLpbrq86oe8HTzhWgYekxETVQUWud+pMc9sWQDl1Aq8MdGomBXOWgpKiw30
jgglFei/qQ9fTnGzCotI9EvjhbeztqS8Drqdo0TpdUMBhhXSJC07gCASajDit4Tm
1y/7uGUfVsWMtK3h1vrDWijbxXAkyt4usylktMYI0UduCdWBEUgKCD0dppfmfpmI
8mEUDH4ecgVMJbHGmm90nfSLxKEC9KeUZ9Pm3PmVyD7ZZgJQtTqBjmAeL2Nu63pV
UoDHZ2LuP1SkYyMCqas5V+tAPpeshUt+cWiC1zdcFaIh2nfnWYMzLtj4XqEDx1iY
vdkYXKc8YCCXzHNjaV4ZUqdekWlnEw3Ds4NGKs9EHp6+YPCvorB+BM0BxlfdjJ1G
AViS/o7w9ZRHxCFv9Yaa/og9NoprvMyEb0rfAax2Ixeir58R9J0H4W5JgRbKMrs+
6htUHsNPIUwq7mRgABANx8LF71PNQJ6Q7IuianVh3eOqgxYwBdGYr4OCg6DCPkzp
6CZAIxOzlodQXzlrEEDc9NxSDkhU32yIRoqdZA8ZVG7agIqmYHhnyQ/qMuZOHjEZ
3cqzz7/TxhIgBHZtkUK7vFq+40qj3WNhZJvB0tiVw8GPJ2S1JbC4wBXUH488zqtp
vdizfDfkLWt6Opkbb2U2pbuvbrJuAprf81iEADdAqu+05WFb4bYttubi4l1i9JVL
TnmSBfTLqZdGGdd9HPqvrmm3DD1jE9fmumjQoRoM+aolSObhilwmTJ7CsvoHe1GF
WxhCeOP0Kv+86gYYWINrDbIHevq9psXnlNHauuSL6j+GntporOx9Jmn7uaCDQVIZ
c8uvpoHlo2DzbTEhOhjpVRZ9jMClN83XKAQXvoro7Ci2QvaDs7a9NVYzg+xKoTD0
jS70ouJBKDahxyG3Ptto7+TbyIHXrhEubDhYfj/FxfHn9pQF2Z+3xC5XwY4OE9l+
RqiStdCBLHDZg5rtQgIdCdiytCYNYORvK3Mfon4Q6hLL/ycG2kXRk+8FzpuMC6Ww
4RX+c0+O1AxZsa6x4212VaTddVFvgtn65BPnsFFINoHa/nlioy/HQMRVUvA6yrG2
k8sfVqgjsT0ri9MJOTcG9X1aTSDrkIr1jBbIGRWouTWWEk3RRySYDJgRSOBl1Pxc
s6hJzQPclV3FQoY4nen47YcAqGv6JK0yNdnX8syO3rpmTmroIlb4pQLP4M2+fCEN
t13o9nQR+iqRV9eU8e1cvMGU7qLbDHk/JFcoBuKDpTKtp4fPAIsCRK1GOYRs3v9X
bMxNZ9KB0pZ8hU2puYIPyYIeQnoKwvVszo+T+FSNNtYL4IM+68VDSUmsfdkmx96+
Dp+GOXvgFrwZMxtjJrW1BrAxKTK3pHm03gb2nsrSoWX0iIdryHNOcLiPT/JECPS+
1967jI2rOmtXOz+pAMJxFJpL7+S4jWnHQfCetfZ//75IjBwRyqyfMiQpHS+sLMH8
SZ9OOGAN78+NexrBtwpZ74PFw5PGFOsTJ+wCxgYCxDFxUx522INQ51L1x4CDAwBs
1IgVmwin4DiXdusS4nbZfjGipcyIN2dlYSdUqMyePPiw3cGdN6gDsdkogVQGaYLj
U0MRhsf2jNaLdPblnk4PQmPfF4IUeX7tyfwbJbEUP+IMwC1wLn1A+w5al2ytGJYO
842LB2YBHInBFS5tdjFI3H8Rne6eH7uELEo/fIz76Ywdwtv55sxJjLAnGPK4YST2
tXXX72+2jHD1XR5H91e0sxQJHarzLhS3IErjAl4tWE7Zeti7YFomFuboV7PS8MW3
Y00kl6ce2E28nSjSErUjzMMi5GjfG2/Ryl+NjTY2HfdtP0XGOSSdkJ32RiBTslv6
HPjE9DN9UKHeyUqF8/mdo/J1+NF19jL3ZIRMvrElvprce8uT1gNiJpqiH7E6YWwe
D8kf5S8EJxi2OLZ/ixEsJRXPEkrPGfdri0z8tuS7SASL8SrdeYbLPYF3rd77DsMd
5VooHCQ6mIu3Dvv43pNkVJnpduJiogH6irMyqCTWtDpliIqXJU4BBo+pn+qEe8og
Fz4W2ftF9UsKdnaIQFlmpZ7WZghK2SNKkUVJV65LADObue1BxqrfN8IrKS6ds+EG
SnAJ902I75r+RQkIhz2YxUPEms+hDua7S2sY2kBFdLuIGhF1lU+6siqgfKcw779e
57J2jhaAGhnOb/rDcyDEjJd9/tRaJbKyV1fmOrSXkmxVMb7KgCvaedT1iIpED4gB
1RjuHbT3GXQCiIpjsW5ZUXTD+MprTtpN5PSSojXwAs41Hj/GAKb7jQceGMbjQDnF
IYTmwpW84ArE5/Y+8YQT+l7liq+OBCrotsXzkdaJwKnqA3VCAiO1rH79zHtiPjmv
R0TpkP2C/cI4JgYbYyPFc60Fqh4g7kijs5zPqPvzypEehWrxuo+lMueeYzCh6UDy
bmnVRUH5n5smR+yReleImnDrOGYuCSASjzSdYc3p47MUpJ+FS8A6z0a+QefWMR2g
o+FdrCaZrfQIQ2sXC6jxBUU96+K1RFCfqmq6aGAHPEvzMgoZkZDu8IaX7/a1jT2Z
74vQzfMhI+wP02enrn/OoHiZ2Obewfs7z2e+/OminBgF1j7Z4qy4KOL4/R+K2F6v
BtdGmdUjWV0LVQJQQoqwaycIvlfhhTdcLjoJsd5ejrjBG9FCGBI0vaLYj1pqDjZu
sAP0dbyWrv1Slm2Co8MNjRdxsJmY69znSWuAIhXz36JBUrPP/nMdHYaVNEZEvyzD
vwJMJO7dbLnI3Jb0m5r/lgBgQLTPVzbJ/FWg78y4MDy/1v2xxCISI//zLYlmhfgF
AdoBkBgAkr46J+VEkWxPcVNQQKv54l6ruVJh6fyOMV7A9yP6BgreAvh3RBHBJWlH
GKa8T5G4gcL/G59NxjAq+LBChhSjgnYM3oQXr1eSzmlUcaZ0kvTXYQ6HkFMZnkK4
cllIVHi+FFpM+VLVRKAKPULHD9WwwkWmO/W/XZU8L75jRyjq1i6rOnvJlx4/4G05
wmDAF5iiT1T23IjwBBWiU+k9nRrmbHnPH5b/wHiKKtQtgvwqWFdtZF0N/lVeoIVm
g2xvsh1OgS22tNxSUt1G985oxkVpD6BBdohkyeaxPrWRJhhw5xJIocy1w3wquESC
pfFcZmpzb90aXU7nRCCYOmDYhGtr3R5Q5wTcjbxCuRDBkA/Sy4b6qCPzOyCC+/fE
O0L5T0/xR4Gv3TtZGy9fZ1XHpwT25FiYSM7+wKHZaoUs3dtzyHmUJQz8ywqjbXcR
os3ctuUgDaROh5sliPdKXAdztvL8aDUZKIOgNPEINSmRztwzqir9EsYjDgXud2GI
9tKje6/WAYSx5/cfJf6+IjKJQ4aKmmbzti1uPQzGOrSMIYPYKy1lhuNEPHFT+SuJ
7jpiP9bjlqR4/Y0LL9Zaw2+uitzWkDjmGgun3GzMm/GCfKerRNoaCChc9ZqTmFRt
W3zMjXa/1QTCRGBuByeY2OXo23CG/glhZN93WUTb/E1KrVygKE4398vVlBoTHzZH
AMx3jSavusaRQuMFTxg7o2pIM78umviJ2gmPd6hDkbrzcQuvcEKeFpzqYCNhHLK7
DynhkbDmKOV9tbxfcHhoLf6+zuyvXB/FFugLDu1mWNjVyJr9Lpam6TXAY9g+tUjf
DCGXVlvs3pnPxJ7OpfXd9tmKFm8tA9VUUwg7G+NPHyHWjAUMqPVIWRwJ3Tv2xdBK
/hzj3Dbh88fqpzCIyMmjuNN+wGGj29KtQe36tIlLpaX+ghT14QIhsHIZPWQJJecj
wx22w5YeaVE4lF+FPuF5sfk7ZgjVZHYokIYjeX6nIcy/5Ihkivu8KJiwLBqy4ra7
IGs3lRP7YZ+Rt/VoKsUJT0810xaaVJv8N3e+wqUscS8fML2bdeN1P0od/GBT9vtp
flmkuBZaCkl1JXHFqzcDzQYCAJnC5biSRCD/SA5CtYxWlyTNiaUvThYB7TrU2sG4
5OD6H7fMqE3KbWh1EHCE/O8OGAUHE4uZ+JUGCldrCLX235t6d3VOzwjvoWrfu5Mv
DSro/8vCuvgapRRH4E2Ac1GHHpWhpMk6rZknXvq4/JPn9IwGLrWibOsm4H2LJq+Y
Tcb6dJqA8O52X0LyU1LW+0NQ0RWocEET8OvHbcHYEF2kdYMHmP6Q6bSeJaJ/PZbe
yqkTqgYPmxnmlZors+SAROE6tFa7BtPe5197BB+JTdaci6DTUt0bcfJKrbT332fk
yoUuVwauKjlGODZTJhyjl2nMOd/3VN0draIWdAq9PUn2gX4kvdcRkY2WsX92eeAB
X0WOMNlxVcFiHhMaKACybI5WHuWgmhlZ9wDeQIzvmTxaeNo+OPzJpy5YCg2iQQc5
PptQM930Ghtq06xksj2/JjSPhEaM8pOouL0ZzWl5XGQZ9GNXYyuq8ZXzlT/VfrvO
0vT45QNiaE8TCydZ+zi9jjYAvKSPvNbSqm7j9HwSUUIjfcQ2PhhMdNlX8raj03D3
/F6TZ9HTt+cqfjOG+A4hW2b5n23BXmsb/W8j5nGyJFvvjjuSgwTNSj5wf3uhApYQ
bCUd8eRuOEXJgYrGhNtDbzCsd1rO2BplKfKGh3LJfUOVsPRu37SaPZM0UMnvt2qG
jGaJEIAAQF/tOHmBvQm0oYi6280Kr9UFCiO4OeQJB3wr4nC0yfpgMv7WyGlZWi/C
7+GCiQXZGfSn95MA+Iuy4p9FwvOIq/ufJpZBvvPKTgtw5I+d0Kpph6WE3xyH01I7
UUk2zcKEyVrhdlmnBc599KDeh5Tw1PUkIldT9J9VT+87INHZ6H27Iw6W6Ai3qzlK
rfe/GbApswhHPagGT9LgYo00cif5JZuva/ekOcQAXEnrEx4hsiIzeApYad3c6pQ0
kwiZtrvf5fD5PM9wIyZD59IZfSQx+RsGE8MMR5AaTbBHx095tIRCDPR1Aw07KEnY
Dd16yvIETr9pb1ces/T6Kn25WO2ZF3O7+lkshW0/yE2fc8nfKS8IchCRiHSYewzm
26pU379zyDgVV3S2QC3bpAQdJmPG89WxY/vV74ZZqzW/x5rkrCodEX9evYgHFXoz
h8i7zBQG3O1MRGZ3riSf4RwuCuaADtukdBR7Q9Mv4WzeAngLeisypKaZDULDk2W0
obq+WVm7Hk4xopvS30WJC2MD6BL8aeLnocysj+PKZRSFPsawQOTSnMLS764Wux4v
i3+ybwSQ0Aia/t2x/R4GRHDIW4o2D0F99w5IgNW2LlNRJDMWEKOeASOgM3x50mBk
3zVVe59XTNTovdKi0zSxs4MtOmVsilTeEg3VTcXvHgL8M6f4uDH+T5eRoktRD2td
o/4TG6baIqG7rp3pT/93DadvoK51Cl1pNlyBciEYl39bdMc4S0waWh8QMsMdmpOO
SGFk8NaN/UTbaFLrFOYBU09HeJTHPd5sB6Z9p+94PocQjQGktoK3c0u0PmglILAt
RVbHcosJjZlBZ7wakidMhDxYTP4zBcxi7twOadM7u1ZO46cojPz6vrvMjOLbM8tG
gyVfLBiBc9KAuO/cEQqZzqL8Fxjwa1sUtZeNDDffN8wU0tz7nQXywv5k5e1oKS7S
8eYuMM+iapl3xvUBrTT5QcOU1EPmm6eA5QZhJG+vOKBnTIgYzUtgBQhzqzLv/gUw
U0wgh3fbyXsXouJJqhmOP0B30sAcq8+PaFrorSvFm6E6mLjjA9G5RzKaCZjWd5JW
GdlxKbXge8Za036xmJFMOfxs8V/L0EdN9hCNjf9Ccx/wV/3yc6fERACEPVgK4XWi
CpLOa9Qs/fAYj6+mSbeIVi91upkCS3vTzRkKUoLi15B8/cutYEdtd84aXBhVHiQV
j6rVRon1yL2Hx6BsVMhNpqo7Wh+NglDefoqvcTSnfGVNO3MzSNfYCpM/5bqOKxqD
l70itlnl0kavFo2mHyRe6CCnLQ9ruR9EXDs3SVDnSmKbyYUGxkvdoo+bc3WANUex
fG8TSJXAqnZafwG4O2+DqTqptnVTcVd5FH0S6+QZ7TIpF/SjxO/qdV+W0HAMfZKk
yJ9P0gH8S4P8usm2kAhhLLvhqK66f8G20B+E8mBut08WywZoLd9UiT3Ugv+0BThr
T/JUBbEBKrHipQom/p1kdYg77bAoTjxJ7K3FQzIQrY7zFOgHGi49RECHRI1z7VQ+
yGJ/cg3/XTnjLjm/QD35Zz39wV9/2J6nljFo6PxxQ0mOD2DxHcLQAWEI4fczJdYD
o4JPzsTxBS2wArCgFOZYCD3nOfqPLfD5sNSzLUXNhcYe1AM75O2lmx3TNa7c5yll
r49/D0BRsIrWVQRoPA+YSg2ssIiV0OmdkeO8wfu9Z+LSFYmCRGjSynFwmOnu0T0r
haxg7LTvR4VoLVmJ4yNJduHlbjF49QS1B+1s1ponLEmptypB49mt9YdktCn/A5YY
R8X1vRI8oPYMTklrNpRWcTUlYJymxYIhm3D5Y2jZfBCI6GWYorwPLKt7CCQy4Z+h
3j48ocxgGCrIipe5N0l97aO9FHBLCRak37b+GAsS2AN65flicPg7FAw+3OqMedCF
9v+4GbQ5KjIWjHPkJnkaFiS+047w/tP+svFPswbRW21PmYeG8DGzB+dLgSiQ8kur
/vf97kG52IsdYsWyvreLAMBsA7LXVknhN4cArYIHPN4OmsmEBaQRmgQ0KHj0BbLd
33o8CglxzRW0PR2XYW6MG4/qFd6guPq121hSn+Mnyi3PdKNFDXftigN66SOMzLUN
I1Kp1NZ7Nn3nH7Ix/OSv/dG+YKcXAcEzInTihPrxlaBztGlfCzjC1uCZ5VqfKktR
qg7UffaQtXpSBXHuKx+vl6A4ruJFWbgfYXocxpGTnmeqr6bFger7z5ZYfO1SWz5Z
45qbfILjnHHZ1DU8x5F2fEeyCONf4yPTY/AYYY6fy7iE8rrEwlSVb9a6vCh0MxRm
/iS6CYPmWYogy89Jv7Ux2Q649Vpw6CcjUfur5qB3E+E8sG+T/NcTpul60aBKWwLz
HrDjamWOHotr8JghCcteub4y3lGpnPg+q0Q7AtM1KnNFDTih6h/Tart9igexjv10
AbI9uvCdnhU2V0L7lOfioLjLgEhKwfXegiUtqM8BcpI/A7tMgrHW48Rd43FraQYP
NVoqBZAAhLjfKoSunMGZ36LC1ko8y5a6675dBVMRinN9Mybmt7tS22lbMgvmpaRp
z9tEGIM4gdRVr9H15cKKyhHUlNlvGVz7gn/x5ScW8fQ4qmEYw635CM9prKVvUzjD
6XX1iJ2u5rC+2791rbe/m7h0cL5Tdl9lR3ZJ940St0fdxebEmshb/w4BQJHQFiBX
ml7wIhLoma+kMvt1eW5nHGOHfuBmTO+QoBeTCHKzyUKQc5OiFSARkwvT1fKivJDa
ZHNrX5nLVNH0jALNXEQzXjF5yO0rJJZ0p1M497KTXsHJhjaw1s2ijOkJAIsiCpjm
DYjbMF1p7OgGntytOjqYff0poJxLMzOogifb1216OqT+FQuRESf9JsEZYAJyAzm+
Opfbgi2unYWrHujB7Z0HCssceBFtqbqBAiO2KFCLESMdfLBsgAhGFjwvRYcPkU9A
Q7t0vu1HBHxsc6dlnr5UxS7KmkNxf1Us0BLXev+4a5y8MingKOQYBzVI5aoTcZxf
Hod4umnBdu4QZuXFxQ5UvnOYc2MKs9CaKPg68lwGWua5q0yjw5vGmV6s0iBU3le7
SlLFlY0PkLrNU1rZiiE/BxVNHuojMhjSNjzhjX30a9piRb4TKn6AoXIrhf02Bhu2
tnY9t60kBO/UPliOC0XVt3Z6Qp8qoRxKAGygmc6fZFBbLvI8VhNrJKvTUzyxXSfh
/84cZcyLwwCNPsPKiA1FKBc70wfwikNPy/Zn5AOOO4BzCmli28gYriyR6hFoGUQj
PgftIRkY4mWWsADM4OqCbY2SM4EIviVJ8oJTLSCzS0exkwiAQ0mkH8DTwx/6k5KQ
cQX6FhGjVhq3Z6HaePT8LFro5z+ZV6tU/RltIeV5Yei3x4Xzw8KyUwAsc2lrRJUT
hfEldTvsC4Nbi+uS+Gyg6Hw6GrgSUNWoM3C7EJq0QA11cs92mmYoswW4y9Y+vH9V
CUgLGtygHcG9M7chIAbuLkofilpuv3Lwl4joGRsxpKbcRjdhVMPqCB3xO5ocweQh
jW4sL6uK1FXK6tLR464m+Da8t4ITECZNQL/9xFHi3obaJb0W8iQ92yhbYjzjNg39
K37WXy3aLUuNk0CnbQPOQHovrcTnLM0AWZc5L2udUoRq1fFI3DcGFAabCXZaCh0V
pWqtQPbWNvbNBrzH5kZ1wCDLtfkJEBlXBWhbdL8sGrkWC709mlrjr5GCRwMcoN+J
7k6QVdCisoRbu8AI4mk1El0tTOXcDBNebKzk2VvjHnRAE8LsQL/uKI/cbpkFMur/
9bdukOjXEyAjGheWb0QU2p2Rsba4dmKUgBJX1AagqGCb/2lA2Tb+TRvw3B7CbZLo
fKz0x81xVSfXT29hqLMBYDvD5EQ/RneYsmDf//2XryzeI4dO5XxBxzu/mFjeABJL
/5Ejcfb4OvDDXM05m2HpHRi2AZ/u9XJLCIZnM2uiENOyg59FdgQA5KOaylT5sICG
MJQZlaZfxnycMDyjoray8VNsavpkqsPHce3TsQBnl5BAxrJpuWWs79QTcUtb8l4u
xf7Cjb1CK/KvQ6DbOX/tmCiubE57d2BCTYRaj0lh0lI6SwHimc90lkmmO6XVBDCQ
OViVDo+TAnXN69WSOhXzhlitjB/9UAEjKaMA8MbsUY4efd0BvVfg/mgilHDWxFTQ
Vg5QtxBMufTwQfdGmpFbZqK9Ta082b8Cvlzl/70RwW0nG4LN8V35YWwxPRvvB+jc
f+dspRNTXUQkQ8zC7202ILIWwu6K32VrOieykRKwMVXokawUbe1wKCj4l5WVlLwM
QUtkLJHkNC/YCMbMbaaNo/dvAqNGZ/3x8ZF0L7bOTndu27Dbn3gWZn9CPh9Zm711
5Tc3qXVn/0xX9Utizz0ZmxmHLh3QxehoGoyQYWbKWP9b206Ona4f6dzDF2V7zxy6
yV2a6b3k70Psj3E84j1+rIJoGNGdfth32cHTqoMbyGwUd5ME1dIakby+kVx0t73d
Mig8XJ5yzwAOZYQtzaf7vNxXyKPjXK0GDJPf+aaQzWg5YRdcUbe5s3pyr8Jhm0c0
YRt33utoBxNOHmDYT+m3sHXew5WoJrsffWLG1dbunDsQ9TqwhIOB//osO7Of+bNh
Jgs7BZs1Z1QTo+ff4xpVBxPUS1wQ84UkUwuufvmsJxCtPIHowuDjegLYSBFxBhFd
jrcRJaXGQ+uNmSPjU6hWNC9Z5UJfd0Hl4KeXZq4R9B3W1d9tnhC8RLRiWk758CKM
Q3Kt+3+pzWExLwQkV6ko5qYqWsDLNfnNn4eocyZsKKECuynXs4ZyCpasOzWFNO5E
r5OiGYgHHxW/hT5t4m5151TEO1eMP0yH7J2ZejbH4blR8r+K+VEa4pe07WFygCOV
r8ZX9/Y6yKDPrNbCSNitENGMRRLtDQ92t0fTBA9NC+XmNET0hoTB+EH/IQ8TvWRF
51tQnbidnzPCtNlW71OWHUDRrENXVbupJ5GLXilUA6ZSOpycc9IqWbei5s80f2zF
297qCp9O1gWQe/+CFlBgsn9AFfdYYna66XNaXdGyiu5CCiWH4m7KdMtgO4XGLXdI
axizfgkYKMXSWkLQDEJzUSgM2ygG619VC95oCWEKb/2eABjgywCfgT8QSxBdetRA
ufv00tHZM6eBcSNSUMl9qNGax8b6169c1XZQiz91JCgZftqucc4+AwxiMr10HgYj
DEDJuSZCA7ehxw7cMBoXumOUak89R05bV5ZCXYjI/K/IwhOvNNTyBMs7LGD1fsLl
8FcOl24t2N2aiS97JYAv7aQ+QAaX9r1oIzNew72sxg4EqHPYgp839LlxNJOUSPBI
KYsH4dFC4BF85Na+D7Wrts469NWdEx3ZXTVTf/+vvuM4UhGC1CgbSJIunHCPgtux
JS3BoZ4Oab+orVOE5oQLTWlZwzPzpojXzLh3KOL3+/IyCp42K93rHJLoziOfqzM9
u1Jueh7dlJ8tom62O/Zzlwc46j6O0G/NXdfkRVcU1lBcrPgU0QD+spGNrvqDOr5B
nEmbUrdA2+7bHwj4t1fsM0AKGArcyXLpipSifYX2O2wpMr1hhG9YXR85boxsOwXP
dQd+nIWh6xCzFZc6/9adL304LxgQoGDCyhSd1lMMuNL0q4jiZp8ylXoIkluCal+r
iaOWQeXcTviuCwE5TNqHOlMe0bE7cUb/JCfDmJzvrdlJMM6N3e+WgQB1pEoSiEYC
+RzNuYtdwgG2jp2oWYKDpmMbi8KPddBHqzzQ3BGMWJTSmouBzMX2/inzQpVFsrYi
LDY2iBzFcpzzhS2VCLHJouWSKegwp6+ZTiLhS8nZZL+S1+9oISm5ghKWg/gWCY41
lFK2GY32VBJIjgxfmw8dMDVNRAomoxNF0NjEhWhQD5iwnwqNkQr8C7rOlii0FNff
07fAp6gMOc/ZzAB0sMWWiIHTZ+BxgnWm8gaMqwERd1hRmDLZ5eGwSkxtIe9D2UCL
UeK2TklTaXhvK5C9XaCmcNJoZFLnNoLGV72zqrz9bFm+HW9OeOWMeqPoHVNh9LC4
39DBk1NOOuYlxTt7nrvuP+Qd+tPlZSrd2Q8pn3bOXWTBeskYbA2q3O9uj9GSeL5V
GUqmcJd8Q9hj1MFUM4S/+pKSi5fR416hKm0OTcmgehEztYcsqME/yfK70MzIsGd9
odJdbJ91vttJWvF4bWw3/uGJMKQWSSFrX8qsKR+5SV7gtCJHuyzSAY3ietdjBPWo
usCrgo4BXAQnvV8WeRD0FcWe7OWOliEctXyXF57iGVje5PFxJrfJd0ew7yAeQHz0
zkAvBK5W6TMwkdlHD7/Tidc5/Jgd6X+gy64HTwSTf/z+dUixflWFRfnIQUWlRy1l
KHZqRsase1CtyGxI0xX79NuVSbrazx1koxjYOo3VlIIwAPjhOBPspK5XPIL2X7QW
qaKiR7PTtMzzlcNzbaXj2XkhVbcimZJpbFg3Vm1p/D5/1zZuicpaED1ybZUrjEgE
GPssI8EY8OE9Rmgz3B1YQq5UK8/PIfZuFCTUFXJ6UTy/rHn48brYdTNoZbHJ1F/w
qYoZ5eWxI4xtjJ8HhSWq8zhKb1U80oZEa7LU+Ntw4OdK8/l/Aul+WXaQRLC7yM9y
6/V656nTWL4w2vsQaQpBX/bREIDO9Fwek1ak0nS6R9vj4Cnjr50zuyEa+uj0PDOZ
3hJRoWtnSxxxSMOQQGmS9eTmdAucJLkjsngO0Po7L+x0UXiadtItOyGVt8/CI7XS
tYU6nYjfIyWl/8g5KnxzKLg+tP7Hh92CvWre1EhJXb8hISN2jsJ15sWvPy0emI7p
fMxG3M9IXfhXvDtr3HvxZzFe7907A+XSUonCbSudmNasgMJFYUZ9CRkq58TqY8Cl
aYa8ciBkxKH/EWdfcNEOkygzY7ZdAleCfIhPH5YT0UkyIlRtttcX5I/ifl3iEm9n
uDkkuHmGVAg+D9YcpFdH5zOdCXJsp0wwekrWC3dk7oME8NtVqdBSF09xMJqrSo9E
HruIYBCIogEMYxmWHbEAIfPYhQrU0kj4FoJv4wKrG4oKlUfc/jaTzSBZWlBaeP2o
Z/QP2dTqf5gH6GiaEXUlyYpGa3LXVNJeMjtyqyCx8KjTuarMdESyOQTI477SGeq/
IKTYWze9skscj1+Eq4I6xbF6v/yP3hR9ef3a8XILWs19ZTiInFBWPgFshL8+uFZt
IHtlNsQPHFsV3K7nusjFS0RpszdEHXb8T14UOyKWVO8iMjYuCF3LXBvObN0OMAEJ
l3u7F21iPH9M11BJBLS8dVpk5YzGVoQ2PDhqhhnvVBt13292EdoXObw0D5D49RiD
Q0/7Uil54z7bB7skZOQQDMhFDHct5JSKkJsgMpKIkN/B1Rn8MS/oPINtOam7Swup
lXuyA3MWFu49gJ21qpahC3dnTvwkfwT8fl8+oxp98RfCkwhVOtbPHssT8z5juEIl
Zn+4w9Kkf6EiOrY1ECPYkKFNssvqlTM6SOFNCPXEhS6gosaO28dB7bZYNhmQpUUx
J+bF7hnHbeQA9BJQYUCKtVnvzd8SNMXqwwVHxST3SDWFxtb/XOm7Z46wTazSjtCt
fPzPU1Aw8a97MzhcSk0CnkTBqfl8RYZhRo0eKnVh1tq3nmav4qvepo0ZNU+gNDo7
ojVuZEckpsj4Zqn9klyNhH7cPq4WdsTOqP+oXCjRKwPFwvo28cTvyAT3M/DM7YlR
o3+/yJ6EAfl54c1fhgjFtz6h9iksbHxyk7m6XMV+bgXcGiTZ8VK/hFPdHnA14iOg
n9aU4J7uFWuGeHO5A93iddhUV5JRrP+iBwOYK21EIjtj3t265mWCk3t9/XQddToW
j/5mlp2iToDU2Hggnbiecu+NyTcDyftbZFmGFa8sy/DpKZT0ChXiZoubaAyMOKUt
gJofW6LPZFQIttWiEqlb4wb4t9cOEWbiLBHk0gY3E7Sk66bHPYgvk2SrTbITdiTt
0clb7DfmOZ6eS33W4MMwEF+TZsJPZjU+nURfvPucA9I8huAKw6boJ4HllrQFEmKz
z063dSu9ekMVRhlEohT1+swBgVDb9EoFwsyC1oH9v0GqNWZWCRdZGaMCP9OOoj//
g3F6epKvJ5vE6cD6s4bAYqUviwvmtLT0wQ54NhZOSHQs+rNGoe0vvCZquQ4rqnhJ
SSGDvIR5NMhBIlCW/pXZbdwhqakDJwlxWA9/ELYoi9cjSF2Y/QBIJ6cUQ5scmUZg
aHNYY+guaHP8HGipVUiQxZa1El5aL3TJTuhhaHpXKpmbYS6jrVw3GC+G+H4MsZv1
eGjMVM6QNllGqEYcCAx9665QhP6s0+D9IaSu+x3mJVRVPQYzr6ELVt2B2pnwCP6S
Ttp/jLWEAif4Cw+Hxa5+orl8HluDaRnd29t/ZBz12B5jvQuEr0UNpS3SitVzqGop
RapjIqH61prFo9eylWzywpUROw9TvoO8GDwVb6BNxqYTGqPBGpP/FI7RZ05i+tmR
yvDNy9OLIcGJyBWnkUB6N8TN1MG0sscIET32BHPC2W6hXLQTM8Iul3J7OhiiCJTS
H6fBw8kAqarUk+0qmfVR9AULEmiD/eenTujvjJvlxdSpROofcWgkHFyX1pAB/A99
8r6qLHTOuR9jvssivMVi2A1ynjcZawtMKFmzY2c000bnk7T6qENGljcY5oH2znVe
c8d4KE+3HSMwr6X1UJKu1qAp+jv6Fim8OO18C2s5BnPTu/ngw9cn0ZigKylx44QS
5hsnMkr15r9WWCikyaEFJAYzEvKM4nyCQJX/ktRSsa4SWYnYnHg2llaJ4VbGXUE9
AzhRN8LZCgORSL2DcJwY/ycdseZY62IIi4C5/HhpkLBh6lbXBH2Glx8N24Ber/F6
CtzNhwx+b9yuyOxAnrgL3X/FY/uWLHpsHcyYT05YAuhxmdee2YjfCuwyOySRDA+b
iOQIzCXZVJ0hOiGk8l1tg2uVdYFTevyt3yrWsV+weaAuCgAoXGryaPdInMGFRyIH
Vg4R0Hhag7GzJp4vZmPqCldAzcNDea0n/BvGN/e7DbXoZ8zbeppiRCOZ3t53dBB1
kHEG91W5xIKBiSNGVvD93aPxmn8XsN4cHB8r3cR+BA8DOZ/c54gtnc2IxbxbjpRF
1Sx6a39XL9CgdOW1beovB/R58mGIYOZ8YrQI0jncjYItHgBi+WFbBu9TJBVbCE5X
lQ0kFlk17k8z66VKTqBBw6YCTNTBfudRxgGFMATKtXmSdMvYVAwtvOu5dG/E3NaE
aSIOfhtHPkx15R08FeHLBt4Ux0qxcb4inpScXag4BARr/mPShH1OOXQ5yyLx2odq
umW5Jbi78W9xgEBCbPHCRF404vSiCa0fycxQHzrhsOpdsYih+LwIjqeVf4OAZIC2
DEk67ND/6eQKPWRM4TXp+iLJisUvSgIJFjvqXC+6FgMacIbbmhhT2j7KuiBNBjiK
XVBsYKUuZLB3qbSYdA4Sz/7NZYxVK5ylMYSgEgiEh9nG0V1gYlznbvsHXaWdDGCh
fGoqc30EkStQHIlQGhqFoGpq6+eJ8p4BPy4mFNElXHJpIzC6pacHvhnSXhXczBuf
2vu/ze6X56d9+eRtc8BJKJqmzBjVkUaJmzItWbhFikGcNphKsTac+JZhEgp2W0+G
+wmBFm4uYXY7rkLRakafoo9fX4bU3nTbOFTVvjkCRtNZzYVRKOCoC6VUgK2OaAG8
kn1TL+q/7fvwgMU2sjwijJgvDYJxhb1drf1Fl8yDF/zePqTextewCi+63DkZtSmL
7neQ/pMTr1Wekerh32bTQNECimvfAP4fRpsYBUMYhFvtRVMjsEd7cceVEynALUrK
kRKlPey9ffvwHZP1ghmdSG+LGILxV3aXw5l9Wwc1oDzKf9LPSu0tEAVS7NzaB/nd
fVwIn9FN8vMT3rtE8IAG2DbEBYf4ETrEY+bgFiJbh1vzunPUglM5TqEHZ/zYo0qF
FMpngj06LlTt6uZ1LKRKAKtuK+KXyooVvKu21FrFBK9K7RnRwqV1z+RK2w2xlC8N
HpDI7V5fvp15OyVjAGBTyCv4IsH/5JheENGWwaj7MZvlQHB7vu0wVkZ5l4bk07CR
nDWHuSWua+doon36QrcIVNJMK8RL8BubS9EdU8+4EfJuxEdhxSdKIKHHdddWN4TD
nBIlE4EiS0JwcKAqSRZVB7Cq+1L/AYqbDPfd4y1kjJFUgoma+nkCaGMB6EVN1T5Z
qE662FnLO8FIX3gzvi0sHf6g/oS54BjDIf7MtPK+gYciTpgkCvu0ofVLyOytbfNm
9NfGq0X2hut/f2E3HPm/9wH1VzTFDIKaiHnRNot7iBu/bq04PqTiZ5X8NpECcezm
Uk++mzv03wT+1ZZJklugBzVh7gn8mZvtBm1IVOJvRlb4slE/T9SD18v4YPOnn2sz
9u+zqV3xStW4gjNtn+cjLp7rCbtlrfNIEBejaYJpsqdzZm5VhRdAwJn0Y+Ix3h1X
x86Ew9dUe5S0L7EbCE4qtjw28STTXW/NU5/e5/lR00xGzea69Ny3M6jzEtMmb4ek
yLEx3WP7mRUVOdNfx/TiHtQCyg2EnzhtFgqopo+i/0tGNpvs7FBjycqcNC8VlHQt
P412wXqooLnVIhwe3r8SXONuUBfo3sA4sEYgjGsaY4SdHcKrLuLeXwddA80Kmc2q
O5yu2BvakYBI7jYenDG3qXHsqXnhwuoWn3BjBNuIx+4ARwi1EYKRK9d1hRnsXZmP
eFMrZ9YikLrw2auZRx9m2lYiD7716c3J6DMtdNbl67sVp5PkcRXeygyP1WLiKwFP
/iqrxQ/WS/8SA39B2jeczP01S965LwyA/hHW/ZoXroIZlMXxkFbDq2JcnbM8Hfej
oDdNMecruv/adzPzAXKK0by/CR8sITrGWD4G9PGIQ1eOQG5+/qYn7ME0jcaCqUs0
cQhvD/Yj0Ulg/2OwQmcNs+95vlI4wR35IPT4M1lHwEBAgLL2jxjWG/v4ohic0eX6
1oGlMfUs+rZ4Y0d5INaUdgzIQcntakmIk0SNGP5Qa8K7OqA6Eo58DJmMbqLIO5FU
8E3u1s0RYQd1IB7/a4iFudbYItSwVZRpfIlTPfeEWpC6zZ+OsHMXjBM9434t8X9G
WJMIs4UtLvc5QpCS1zpTFTk7YFQe4mbnIVGV6SURJ+9FAhzU+Q3TK1pn6IFALKzj
Yozc38n5lTR0M4GKetet0XB4IouXxOWhreT51EQcw78lO5cWIc3u/sahh3XQIl/0
FpZcIrq/+4fpyPty8abAJvCfbX5dplxtVq0G6IJVfEOfwiogmEr+fvEui7inTlwz
6pBfviylQv1Lo+gjG9BUdhsLeTlilNvK5NsXozbiVUM0PUzqwqgjPLPq4CuDlHo9
av7ggxkAmJ3CxjeL3NIszJ74OqWGl4wGyxHQ6+dLbvizTHDmtJiL0OI2m5TX+U9C
xbW+qCMlbZAOUUjkvr8YxPW7E2FnCOgEa7chCxSs3RGZhi3mEtD8HiRbh6OMCf1Y
Q3E/bFCpfcH9yYvROOSLKU/hJYhOjL/2DDaA/AXJf01eloidtQrXeS4s1nxhYNrI
Ss8mDCmMJFJTTIcKwzUBGldiBqvCWo8wfIvIp/vXs46nlh5XVrOJamfYElsBnDpr
MvOLlbCw/pRCNX3UDIpzjdDfzkkjUldsucPdmwdyrKsDVoPnDPmhtHuSMDFH56jV
X36j/yZHdscsikSgYcYFApOIqDfUorPZegqDrMrqkxhnI/vs4ql/FxX6kphDBrB9
GSW25ynEZZttKN1dQBdaDy2RCwSUcCXj5Njd2TuNZwqg/z19TwcjlWJy4JGgSHUv
QZJ9gp8awpfcabCrGHcXCg8fTHdROAqrWFyJXPIfopNPdv2Aefbu4GpaVENKM91I
ReUV/wJQrwu4VOCCUFWyHVwoRVb6mvCDIyU28hnNnl0bYixvRJFCqSOPm8b8b4rO
bkbVKv1zha9q+VwNk5/iuHbqhZ16e/WocMEF3Fw8zq6USd20/VeIJW5Pu+rfiYMa
UKa+KSRDzL6u1Ygz05Z3yMru8pgoJYb5UKE5zObGND96+7kR1BQL4PWhvppaoPVi
nHZiSGHKInfqBdxwQHglTG9tHEFz2+vrhSwc2AtCnLz+k0e1zWP9usCWEFpbOrKQ
mo9nwShX6wVSec23OBgeMG/oluO4+Xg2fH8Qc63qxiATcLMgc+q5Gcdxln9FgIxW
vyNUu32lvLVkvH0f+i59Ouhj8S2Q0noU2K31GdyUYmvF0DaoibswNwyW/GsQDo9I
Yi+NPpAof31tqar4VBMjIjXLCoeXOpzcDtRlNwtbh19Q/XRLgXCQFufIxtJAuGWa
QeqJbTm20HdWQMoGTaOUSdIN6Ic8ZWd5F8VL0H6FgudsGmkejYUTZRlsEt+pMmX1
pyuuNZscKG7dXY1CuSJwqJIwDy2HJFrOy3wqdEoIIL31k25A/67UV0Fv8WOPRgIr
+FBoMP2HucrJBLW3VikGs/Owv3tGw/8SqHepwuM6HMEdv5WIgp7shyLXy0KUZ2SQ
n7Thg6h3wl97c0ptp1uU9PU5e0GRBiO3l9TxPxiI5TqjNJzfhK7S0aNKdFwL96XH
IkdNWpCcj/2UkRNZbSb+DBmXgu70XMvwfwgCRjW9OuOORsCXYHh678FbT43BP8tw
hwjHcPYxZUoyGu++R8aopCXeYXl2k1bDZyhEl6If7BfqGY46EIvE9Jrrpsay3H6e
/8s+Jr3w4N6teTrgbOZHlcfteqFxMOHP6Ta6hsy+HfZaXhAPRXUHbdHWLYwhI0vr
0xMxeh6IeVOxobpxaC03fcVOuAQGP64sPpGkLvRnrR1hBPHTUmqeTZCfE5wG5Rz6
f3CyRRn3/oyt+fGpeeqHehW7Q5fsfa4PaEOoTiInKfYz5bM1fNI9t90BMBmtP/RM
O4qHi0MtzZIqstwcuSDi+qoUyU3IyBLv4gGR1ihAtQndW+/YjehAlGbg2LNWODpX
DGwcfsHXcfjc+/jqnH1/r1Yz3SXIVt/UU1H/WY9LedQvum5D4Pp4NnZu47B2DHcP
Qaewic0gtndPtXQ/DVEYAMZgZ9iYm3UiIH1iMX2qG38L/cSHNuFf/heUZctSyV9s
vEsyQgRTb45+f9nE2V9GoDU7XYpcu1y+6sXHORdRi6C9xYzqdvRV+ciWhQok7/F/
hjohD8jhnVPxsBRwUmk1GmDh6ccyo2PKIezNm9vk81F6DuBOedMqNLm0TshVWNtI
jcE+B+0IpmWXV2OKOHm2KiHti73GQsTI29f8Lvey9o3bxcNVljJ2RUVRpvamr1Gl
tTp88QWEsosFsJnGSSJ/sOWIokgalaYMPPQ9xHGTdPyJerrTnYARSc4d6nvZyB2B
6FjErRuhNVChxL46q0ywr0hI72VxrYhg4MN4QI1Ut8STF6vDXuQPMEJ/g8u/vHot
YrRsF0vTrm/brTcGSZp18LKCGc5Hh1h2rkESFjjaoqcFXEwsOTQ2ZUBdmv7+r62K
6+UwflLPsKroTAcrOpX6e/1RB4ENoEvjb6sbvkWh9BL76QHK6mn92aEh2pG7Bq0k
aM8pYdwzFnM8UeO2wvxFxPEfMO3DtcV3iTLmgOwF65djewExGPDWQIUzjSW5FaoY
ml9QQ0TUCI9+97dcpCYp0nyBJQMU3ACdTauRJMnUMEwbPzxv+Q3gA62zdRS0Hhbp
sXIHRgLCtPuJRPaM1M+BGYNpqAyf26UAE1xpOrFJh/NtyksHvli4IVGc4cKTo2cg
PJlPqidBdVYYvb9xvd/NIfvNegaTZvnmz+bxBIv1lgxkSrQ2G9UKU+rmlk0x5WDX
IGcyVLsUzOtGi44SyJr8Ywh2XtENx9OWB3DFzb9b6hr5gRe9wctGuQj849xkcmT7
fd0gRknzkgDqdwKOt/bDgiZVh93uaKFxUD4O5N7KSW6eZpGa7cFE2lOwYTodncLh
QhT4W4Bas39yl5HvjV8kwNxTAFmCTAbb1zg7rhw1aZP6ngqzc3RYeS2/EDXSZs7x
KZPbjU+wPArRRV+OFklmiKvbw4Fmr0r2wzFaxUMzLEGTe0OwwMlFtRs6uY0V7u7T
eEOQgOgimUWD7x6fWqTtWTy6LfN/lydipXg6Ak5NqDkIg+EwnGvgt5vwKJeV6iAB
qSLGG7deAyxL4LEXVOj1kvsHPXO1ZLoMLoJb80z79MgZxQpFO141Z/Iu1X/XjD+p
3DWFUf0ZVl92iGQLAOoQyRwuxx0VKz/fzkYPY0HTkLQvblI/8BxlPqv+7tRLjRyp
b8/+g2KoXuOqL7khFBHdtscWDLR0+uvEtoP50W/AdbGViP8OdAmA0UoGtPtpW/i8
BaLPcmjpAucyt4Dp9Bw3L3o/A64QerH2Ik4MBOD0A0PedyjcM2hQvJyhCsesO9aR
010dcEt8BwpnZkVTn0y4SWJ7wyGg+G/0Hc77tN6qhSZgwsQzZUkS7l71reJMzPb3
h7FQMhvCGCXTLW7SHy1FV0SJEQU3oqb+pS4xK0bqsZY66+UKJahoQccPIWoJKvZ0
CwiiQnydyY1f3Jn0E1/h69ikN8wcbjVmUNhlEs41XRqDyoMXBbtTcQltmh8EhAQy
Bp5XEQqv4Jvz8FIUx9DRCdm3y46PXIj+VarX7bKUbFmfHrmythPIIpQLchBbKig3
4zEiPrx8/yzvRmcuughcUhxMN6TI8me9xNK1uqRib9f6BfwaTJVbb44gEjHS7hJ9
mTFiv7W/nnLeId3T9RMuZWQpuwgA21ossVdJJp0w9MSpzSxLoEbh9GxVaId1imOV
JCXyrrsIu9FRsIz6CV6lxz8Xwa/tD5RcfxTwvqdUn1GSz06PYoSLUCzsH4WhQcvx
8f86E9oQN3m+L7cqQuSaIZ76rO3KXGZhVwIbvfuhQbQrmPKPeV4dn0Mj7gCPg7dC
++kd76n5H8RvCkKtrMaTBtJtiiH39EAwfAU3bFJxAof7OTfBlNuBJLLdRmnFUqG9
5PmrfjCftZE445e0+pRS9Y/tjNOl8iSxyZqBe6F1BP5ZtKsWLjEyCtRmmJjlsQZ/
TYyJkxRhRT5gkAWYYHgLXM/hXVLKmH1DlyVMPUTd8aQG2Xkjw4GQuunIvEchI2Ha
D/rol9CEaeIs0F4VNXZhf2D0tglkR7X200+TxtiYwxv49pYc0ZEOtg7X6cU2JOCK
nqWW/663GOEyaRlDhiwgs4chK1hBJGvizL2xGmVcFbUrc4It4z0Esnr1umZj54Ih
CkLhoQo0sKZzfBaXtqy8i6NES8/9yopZ9+UFQqLZP+/7hJGMOhfzgY7or/dTk1o/
Xc8lHiKqM3YoeNBp6kAEO2KOANsHulScaQEtDXe+9Rhyrn8CRwIctV7MUkArIdc0
9GOH0mDRO6y4UsRhMeEo8k7NXisy+sfcNfXyXLAVFHgvJf4Pk4lG6w6Bt6J4zrPT
p20TOHQg57riBj7VoVuuec3LOeX/qCMMkkhy6F2TrHBr7EkIY0DLGU1KcdOL3TPT
aI5UEnAPDorIfyo/6BS06giWfKPr/dGkrKfEhtuBL8PNPWbjd4wpgmQ8c1nWtH1c
rPIA4O78svbeX/t5EAoI0essH4L0pqEKbQJcsQVcw5OigWyEDHCPlbDVcZguxbdS
P/CvYmaQRNilc7aIxw6p8hQWiCEzJG2opX0J7bN5BvLFUNvScQCt2KjdloSl+Pxe
K7Cp5pwLCj5Mdzrsov8HjPqZJii67IVQR4VCIjgvyhAp6LZ0z65sZwr5khwZEjgD
0Qa2olUy0BsIDaWM0BiYJhQjOfr4pZOXhGvVDK1CLjpUM2R4Csf9mFYIMzB8qx1O
E9qA1uua+x7a/ol1DZ753fzVNh5NysdrElYR02u0mAZMpeXV2HbBZ8B9qoVsYCPZ
be32Qw2nDS9I6BbeQ5y8kjUhEL2vdrqUAlrzpk5EU+52QIH2ro8szu8/fzNYNMxs
GsTstsZDteAlSWGa3rjdYMAahWJHLLiercedV3/VZ/ZoR65a4uuX3zEizXgbjnvv
CzLprDSXtwxNuMjS0mgNkFUD+aqVDNyl7zbdUvryAzk1aAW+Z9gWi1pjwcRg5p3W
M23z4GbqAlhmEVbMDdrshiizObOUmkYZixLpmmabNxWjQj8qHO2IzlVyd7uzMBeM
ZGOO1kaRFzt3ty4ZXEpT9UPOYne+clnVOUYppKZL8J1/y/dr9Eg8OUU34UPL87LA
0NSAGAQNDG1tqHgOTebYVdw064IImzXQb7vwcs+ZAeOEMri3Hr0ogax/En2+X+BO
ez3n/vF4IzYjtjsnmoqre6JfrUkdXHV383JSbS5+1RQGopwg7wuHhprpp840UgJW
0MmRwouVLgeGxexRMleUIS+I3ne/IVY8tVIP/p1UrBHKChc2Q5rLCYtd5/JLI/u5
rUObJnhoTMKaWHXqhmF18KsaFKQGs0/zWj4XFr6hWDsF3dgD9jH1KKtIgEKCWTRr
sQeRKVq8IBiJ/H7zq1JL9GJLtEMosiKqh0+uGCuC+Aauehec3a89D7yV60tJs9j3
znR2VKZALulePVjZ66phoHGKji/Na0jEZjRh6d9V/+EY0LtmWWwGy5BdRLNV6SQK
0jHhy9vxNrTOR2cedGdb8uUph0+7cRk/X8AS+Bgh7m0xds1do9sMDKL4OYHr3Zng
uXxay7vkI3mStpD22pAOWVqUYwutkrWivu+PsgIsK6mhRZV6zBHehYI8zWtC+Fkn
E0CnrH0i6PSmAjxliPj379P90120Ynz6UtRtsdA4ipsq1Codvuhu3wsS6insmlTC
UKtGVraSJ5caP7YRzzoCWcwRWjiJoGyERG4hQO7sZFYyIHLoCaaCl4roX/HQI5Di
ki5G66YLThdGdUaR+3Ve/tjT7hFFGAf75/0eSlnXDmgsxeC7LYHyGIfFvNj+1jQR
ffALN6rjS5N9UlcmvjJYMH+O/ej7Dt9XyA4cu2YDborf1FyfP3QL6i/4WgcnBkuA
xAZ1N1aNzkCnij+kpm4UxqL4giHl3zgQUsupV/0/qeM0iJkMU47dJsC0FklkzUZE
5FCzTBUtAFAVGIajulrnV1vd54YBFXSBHPzbAGQuJKGAYy3OgMD4xygl7RjFSRD7
6RvWSb6VAOMbU+7mTjuZvNEt8gvvQqgRTu3bhvgcEC6YHxRYOk3eanHNgXf23qIn
AxFCxE+Peo1ohhr1FIUZzINJZKHsNbJuPfljqdjVFVK9bBCn1ddcOA9xs+91VSjf
dqZ4MoThsfiPh3OfUP3uouWNAIdWjh/RA9lD+Fs+tLlBVWvbE+arh6jhSkUsb5zM
Pg7ebaezAiHdanEWK+KkdCqM3v++pbY+Nbz7Gfw0JWFa0rVXpZ58v+aeIfrvZqC9
U6Uggmu3m47g4uqzL7nrU3QV9xqeNPiX8AYupft8bVmRnNYvr9wGIRTBXNAtZZ1n
mcgxD+ytUUgk9so4lDOXI7cJuqPCTuNa9+nPAA3IJioaaqep+HNUmjpPYoj6/prf
KpeNtipLQKxBwVYpnEZal4WQUHnnZ4kEgOLWszLaJMvNQNqEsNjMUumgDIA3/X6D
kHxKQJZ3PzEh1SWgogZ7ekL6qC/N/VqLX4awFTAVWrSNFq7yH9xEfaY9qSIOaOaT
Fhk+zKt+14/99Bn7W41jMmzd+6pTYB8fVb3CrCFZHv25Uh3QMHnJRAvxZbr4L/fw
gnN+z71eh3pa16HCQrxtccBD6k5NiRG6vHBfkJEYyElfYpq04n820UhvquHSTaaI
75Qp/fGdUmmQ5VfF9k4MH4vTzV+P9O+FjRPxSu3cLVtnS3mQZNaeB1sf92n8sHUZ
fPxCMg2AB1EZ1AKfTSbe6NKHD71g+ZLaMDk24aD7dTC75OAVK6tNrE/QhoIu0paX
RjOotyMHnnqUl3SyiruzApiy4OgwaEDJBvTaOXjOO+Cvo0P6A9Uck6AKcYng690i
vwAFjbUVcY0WVt0VgZ5SvM2IJXDE2/57/fnuVS9cAi/ByWqKqmeVd9w3RvQijhp4
wK7qpAfctGanUKjJUT8SUuU/+jzazkgNHC34pW90DG4mYbXqrp4xzkiKEot/8jtu
mqdA0ZSreMrS59m9WjB4f1EZDkdg4Mm6hgUf8oVoDF3C+8LOlvrfDoNnfJO5h2WJ
MXO1ZEMhItCWl/7wNQQJCAox8u44l9guHeUi9MKL1gjXgm/+K40teuF6fBmgu2PX
Kbr3L+ckVU8A2r1huYi70Mox61wCVe3y7o/9Ncn1/9hs1Ia2wVWuP4Ji8yjHBXFP
1iASqn5J0yw8HUeFykBm/OEJAOSiDX6shYI+DMsi2TmoghiE5v0M8BaDW/YgJn1W
5dT+E57iN8h3ClX+BgX0z068JXNghrWT8SUR8j04PbaLUhsU7LEAOuKIFIKMkgGI
+egRHoErqH5tuxwh6YyPpoDOz/kkPviJZIAY2vNtBHWjWcUU4UrM8MU21+VGoV7y
fZwRlltqMN6FX8FIy/RdXyMxC2nq6duHHlfBoha0KvEKXHRWdEOssK9kkT8im9rH
RVDQ0+JFn7vWpFOnJoEKjGDJkmhwDdj6wCZbW8/oWoI7MaaARmo2TvlYnyn3Xmw5
UmR870UDTxrwi9Y1XBNjMoJQb+Ftr6l62Jbn1ubvkM0+8TchXkho9TIT/r94VEwQ
w3BGPSbtcvLLajBf6YM/YMvyFeOxbmtl32zXv2/8JlHynNOotXkc3XQ7BE+O+7mw
OOt1r8DZIeoGslT15VoCPlUPFePCGe6DObjzAV3Q0dzaIL2gp8wxhRx/mNTekGOF
B+jr8kXxkbnbdgd5hhKtx6gODf9RFaw0vVedrfdEudpWRmGP7T9ktL0oMQ6frYPZ
D0SwuGUa3+OiIIapNz9IHM+aEIPV3AYnrVLvFstAUC5A3fiLTeS/DFMn1eUIABK+
tUYNi9pRmGR+VCT7LHQDng8AK+6sSxxJfi/Km2k1vljcGe8MbN7dbvFIX+ROILvj
PuHf23EFK2a2sk3xtREbrPIBV6OQ3r0qyoJHyjqO5BP1/w/mjGXKfVLjdykYfJYz
jSPuSxm1GMK3Hl7wWHzrgdrgti0QsSHWfhW4qfTbT2L/LFyzlPzU4BbPG0vhlgcl
VKfG7t9jb2x8MwZVxi+Jwa9XSDkmqVggnomv4nICBtg2MClQmShIy8aMnqk4izch
+wTvgv1CxfTTYas9R0d/n2FuqPk3iHTnb9s7l/QNUEJoCZKgT2mKCQrJShUnLE2q
+78HcrZ3kDf2ktJG3o5t0+DMzIpBqHP0yTH245pJgonK+cuee7Bqqnyid+1f+RqT
xPaf455mlPoUuvamCz7QDp7KJoa08fjoRHOTVYslTstvfTeINu2fGnKAmLi9PqWi
KjLn7wa5SO7scm+M9/1HvPGQuWOxkm+Ihka/1z4XQAVq8jLfmPRhpbl+NMBaRtng
lxtkwY26McLaQEWqQS/s3QJFNrs1tCz+TJvmoTcy5m8hY6/q9LYfXX1OrWePEoKQ
4ZUb7h753FTpkclKc8QocQHQdqDqkbiOia3OtwbbW53HJyBGCpDNBoW1xp846jGz
Wi2ReNwN4mQTXmJ/tPIoMuaPvgar4MGkNNIdClH47GT/cYQVqX2mKKza/e9jV1oS
bL/4y2PUyZuQqjs+0tMSfK8WDaVXSTxJgkkwsLufE4cU544BpBUHmlJiKKfDqLRX
ijmlrMEqwHbzId6+jFBMCE97zlYJwnt/wE9/Jug+UcKY9rrJk3sQyCoWnsMYkCbe
B6qoYjJ2HTbNftIpd4y8L+tvBkhfCmndkMGVm0nZJAF1mVyAwZqpprIWIamEuu0A
BFR9EYTywQQ+40gMy6wY9ts84EyYsM2zM5KlhOLZKk2xYQ1cjAjkVfUjCeFQOfrW
77WnRlwoQoqglXBrKDtbsBs++gzyDyl8HlCgy+xjxKjYE8QJWIeXP29xuH+co9Ty
qOz66Y+6VjdZWuuqmZqp5W5GQQTY0ZF+8+mXJ/Ysgk7QTeu4RlHzD1se7/01b19F
Q7FfmU27W5ucMbpeSpVPiJxf/tvs2nncaVI9t3u+zXdW8HhivRyMVX5dC00Ao709
41d7ns7F0ligWv/t6lPTHgRfclbJmUhVRAwTF8PTOVAXIciPKuqqY2mWwY2M9uU5
Gaf9z4cAxJVrF83q+FLWZZv0PExYmOhb0C7al8ikkagG/7pLc4hInyyWJ+KrknIM
ZJaxzkEy7xbgdUP6+IhWC2/fZhLEeNVl2ZMk7Dbnu//nXge38lhWAJFMah67fOE4
lMZxYDsFh9ItN7tpeAL1hlqc0giq22kUjDTZ4vmEnlwm5EYmnuFYezcA+ne/fN1Y
UNxkxKFsEk8mCC/pIYDEyoB0rnrQVpvgcASar9S5XjArtQofRSh+mKbiyuq0UzjA
a9DyhOGokUSsjLNhxyCYEaonIbQadHFCeQtN4bY28sh2za/GYT1dZ86Lg4peBQN6
YzY3VS1FX9/NUEYQJfQXB61fOBslxL/yc1qk/G+QxgA1R69cgea9rnNpbfHB5hFC
TMSnUqeJgFHJ+UR/Q0NT/KtWZy8Vk3iPuttU8H9norY2Cznoy9UEwqy/Mjf4+jHT
GVGMayk2C4OgosEOjtWqsGq+2jvOsMwtqub5F+WJJXn1IbRMiOshz8hoXy7Ld/d0
oHw3nBwL5LF2iOMEkUIJcDgbnhddEzkWa8lXMY1TPCHQi8K2EAh3u/1h12NYN5VH
rkVZRI5xc5niYIsCj+OMEEbQNzazEn6lZNRF4Rd8htaAOzDEcWT6aOE8xuU25q6z
6ZEGA1CBIxWFK2WtryQXfE0Hv9eXYMcGtWPMwPpIypCMM6ulauz9byvBVZN+tok6
pY43K3mqoeKbb22iLtUIgTeeuytbAGEElwdi/1NpLd9qbcKak28Yvi/fMYirtDFT
6RbXc85xaUB3XyK4DamJghMrVrR7l/R+Wp39Acl3LqyrpcuGZ1N9oSFJpgdrXfSu
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mzR+lW79mTIrsJk0RM+hcNwX+NyoZaNVxA9UVrpddfT+O3bs9jbyT0rbGtwn6dGM
GXJp+TTytdtWaBuAnwxOowEH1APIOtIvGA+nwVUnw+YlOnOzDgghpzSi+64M440g
CLlvEy4aUf3gJpFRQROh66JAmq3t1ra4UBCZ2xcofVk8In2iF6+jMcsEFTxHRi/+
nP93ae1C5UMfN0QSa4s2clQMsBnRsiQBHf1b61UXJ8YFyNfI3Sde7jMb8cMZhRHM
yTxYqqm2ILJqNBsaHjduU1ZpEWHBmfj9uGPnzUTpQymTpYrIOWuAhy9eo3mAsCKy
fgRQ1iVC0TR8UvX/8mhUyA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10032 )
`pragma protect data_block
Sc/o70/y3dbFmptIDncEcc+WTabKRLet8ILWi65u0YF7tERyQ4oXjncaWb6EIChF
GosTgPjAFFREMH8qdkYF2C3j8uVYYwLk1e6jx2JHea81C4yNfIVXNW8Wan32Ri/7
3bom7rpklALZQjpeEsLoGLM4IliLv7s+h3eSR1rpQ6hkQwGGFqDmtjXHkWFmy0YA
7Bmyh2opevr2NnetXLVdPReFQ6ynamTGXJv89LAqe+o0SN+LiKRZzWPemuYX3Nr1
SgrIpFc+jcudfhnJlI/vkS8EKsd/1XNPS1cfOxCiqWinsrP2bAPu5ggQzJ4czlyE
PAGJCbHFeZdCMSjhH7yHFUZwS8NctWEnrrmrSf9pUve2TOdMJNCJkEac2rC7dNhN
0GBf7BitMbsVecXEkwEfDhjfWmquC0gEGGu+Gr1ltda+ty4koSDqV2tvXwtrYRM4
xZnwkeEAR/oO8eWXArfZ5B7a7gqoHrVTD23QurN5S2lHLu6CXIbgh2OzfB0TDzd+
0EUPWOtXmbFXSs09ap1B4NI3H8b8S4giv31eL5zUOuQDicESl+5YIWlvxJlqy419
0HrURWtjPeFo2BSKXsp+z/ePj5h8Qqo7CjGb+S+7GEFid8640ShbICLRmd4RfL/H
vW5Ozg6ky+FjoKgxWCkPWgZtCd4FC1r/MupDSzI1JD3QTpd9NvSrXkpmWJNzIS9E
/WNZ/lF5QEQ64HnwYOzHFaeX5mqsByquT26geinIQAjDr9SB0N+mrbv9f0u/blgg
yQr+s8Lmb88FjwagBYOZ+vBHHn2SokJb3isHGVpQlQxu6DC56UOt3kWIaP8nknk8
xZUcH0wKs+xqUoThGnNe+8ePX0O/AhdncUv1Xw2WLKDDPo/KkJBOgpN7qer+1Ga0
0zN3H4SnFUKIfnXkP8rhCnqAHvjz9abC5PYfrTHjl8ym8A0yewQS4yMHrGG5Sfgd
Q3xfj4XDu78/igtWlFV8dHa8GD2YhloQ0FXvz0nr+ogfjhEOsSePWYBOBpmSd8wO
oeVPQNbEKl0twjiCx0QhzX4B0jvHb4t5fiyMES1Nj0OLH7RQKMf0tdAdSU+VNxsa
0yBPxul3GCKPewBVCVgZ+5U0fPQwuMenLevWilzNFTZ5nq/ksMFI+TTjC16vtjQB
qLjNzn2FNe3cfvl+vLDsjiroiMfAIOBnuUmafo6DiH0GJ/kIa7YC2sK8G+P0bC/z
7HjZ5h8db+S7Bplhs6IaVhxh2Zg7qPDcIfdMFA6ptDAQzIhse2joT/ija2tZioXg
d+wLnhaDnchp9r50LidnQRdFAbOxx1HA+Pxn1101U4uqJ730pDneQin81NcabujR
klCGagNhIi34D46HexWKGtJ2unA7yqw0Wd1pfw+DOwQpJCmjNauM0mrdhwMVFbwu
0WJZrxQ9zysD+J8PN8EyLD8/Y3cQyg00+P594fYwNROxDDdLNb/BbraY+8CgC+F8
1atJbWZhV/NhHnKpjn9aZQXy3cfY4a3ByaV+AyAQoryYXUlLQdYudwcTWd0wWfXt
SBqftGIvKZa3d0CG1CQBAsUdIMP5XUotTnmYU6ntNX0Sn2FNWEH63nRfiHzlJvvW
065L1Eb9AL51Sb7t+x2aG60WGDKLMOu0XxhJZ9fUUYGq5ari+uY5/y954Xt7x8c/
NngBpZYRnujRqLKe4L4ciIYsZ0bBmKuCIcM+QbhxlFtKrte+OMN5pLxgN98FuYfs
t1pV5Khj10BsYh9icoV2i1XX/j39UAgaA5FrSN6spiajffOxg7o81Yryb0HokZ/a
1ybIB3mpnwvXs33wlpTCe6QObXLuK7Jpy/yKwP1WaeUND/ZgVw9uPngx18R+v8H5
c/MFQU7AWfsbv4upF2rM5fzy2bR2uNcYJ4DkGI+Cs3oWFgViq3RP22bPc2llwkvq
s63MCMMhjVGIe9dQvNcsvrGo8XtJuKQS4PBPNigTtVcrhFwlCQKdhZgKgA/E1lDY
KPlulwpEtQngfD9m/rkXczN71jOmF8UVgWBUlsUsCvvBksQDd0qvwqv284n572li
kYWyxs1JROuCL/m4w0lYr8DsjZi+xV75PWMAJmeABC6e3YzNill7qmoW50KgkKeH
tQqqFtiM3pL7oVS3ttEdJoEfyy+AihrUMgqZnwbtL4auNIBxTNfsas24d81EQy0/
7kUsMYvpTpuy77G8TjyVtqEbJwotwRAc79kD8kTU9US/zNLysFx2+hmXd8dhVq8J
rT0cqjK1sUkXtttddPraTy6t42NC+F6D9v6AElSW5i3Qdx8vAi+MGgXQPlYEjebp
0QD/kO8vTKTUxAQgMXT8kWMzTmcRSxg4jDpDxi+9l1IdnW/zGuCf+ue1vt80seML
Be+lyIULp9EcCNPqjDguYZXLoo6MUxFAAAZDshZJ/73LfjfsCZAriXSiY4hHV6Qk
6LtpVYgNzlLsbdHkhX/IupKujKHNTWlytBe5nJZdZ1vF8eid6iBuOscDKtAZxhsM
yHcxcSr1Y7IC050cSElhaCRdk3eYm9gQWsahCzeqWLMvgjlA6xZ5zrf5//X+j4d4
RpiUQm6bljtIo6YPifBYubj6QnMjeYpQV9HVQDVBm4j+ASgozI4jttZ6+zWn80qy
pbkcYvFNL9iluq75iU39aoOmDFkQyGYNAofn8TR36Dc+32Vwj+tUZsqxzvrISpsx
/FFkhmLhrV3nJ83P/uvA2f4f9rCqZ/sETdIQOdOcgclM41bCmXr9ECM2jh7oasBN
f3HeKll7+7B7H1dzuaYIpxDehXQ7eSKIs4qzTdn0VxzCQHHk4vZN/dtTZ6tfkwEQ
+N98jyzgC5E5vgLDmFYEvgLs0Ofx294NlVsi2IYKtV8nKTAn7qWRNIjzurmIOSHx
2yNrTJALgz5ryKfTDoNrULKC3zpI9T2WGHuwh3kP93xkw5Qp6KTZ0tAU2l2+x+5I
3+bQfUN3uk25OsX4NBmO5uHxH1F5ChTVMtzPF98NPE4vMCKwOfPSuTS09dTwmsNq
2s3kfHmrDbyPva1P99hPfFjGyP5IZFkYFTlOEeQCxzOOSJed676jTA0JT31oszLm
r3HdfVQBA1KY/UFbX3OOdS9IBdQJhIA94ocnf8cdIzw/mUDiE9gd15ieP2ABIxrI
1yzqkRVSwEESi2g0wxrhxDgt7gOfxYW4q79jEHrm5FVfrv1aGUrBwhyiAVACSULX
uvwlj2USP/+4wgMckTy6d8keDeUG1QbsuAABTAdIwnNCYIcyaq8mYk8amQ1hjVqk
uxwfgRjQ6Vd/BD1kRLCOhyH/nFkmBe7LMGCSggFTM1u93DWGZ2p9Y8b4MY5HCwjX
t7C41qITlYwbd5kQ//WOW8uTdIvYFuDQj9wdOrLaUQHmrCxc4c5uPH5AJB00hBsa
KDwlXhmDOPqmHsCy9vsLT2y8aah1NppIPn3VoZn6vU43F2OozKdLrIY29XLMNRXU
zfYBcbmoEnBLOfkM2RxojMdqvW6vUjsAw0u4zl1B2STtLBx7TCg17a7LbWL7ipgR
QVDeiyU63l5OZdH5WNVJLvTxkZ6seY+PPjBW/J4S56gim1xwYzVgcBhNcTGBaflw
BfQhOozNkB1re4KeaQo1frgMXhJLK5qgy9/YPZLEa/kSgnygqTGEFZLPS69bH1RT
7VEexKaMvIb+exJ3QKZzz0cfmEQGZ2TeiZ4LL/thmyc62jLPjbGEw8mZqFGces9x
VxhqiAXc4XBFvl5kAyTUSyAcaNwCO+8fQf7wxcJPdMJ2HcKMKrfDCQduyU1QCObP
lEDe2QrehzbGPK78wHj5kcppbvGrViW+yJNDEQAeA+UmyrWtcDbIksdQ4q/dW4GS
FDIcoGOG7QO4vH7EzTPK32X4G/oxbvlLyroajOThH0Rn0Mmk+61pSV8PAH334D66
tZtaNOTodavx9v7y+gJXCGSesJJiHrhBgA2VNdhzwEhBQyMfb0HWvZ385FAhDV9a
nxxFXwZt8J2H0Mn4MnWhuuXHd59owr3wz5/kcKRMgh3lR0f/bmYSGpLHrWDy+2Sz
jG3tvBo9iDbjN2YmtdVFmLqj7anBBQuk47y2Y17GMlRODfwxV3IWJLYSlT8Fy4JU
q+Q9TYyq82HuWj+wkF/ZQBQfsWqMxA19ho/xU4aENLcl7Uiq2JgMJobsEjjQf74T
Z0XpEzmOoYwGTJAl43V5xGM5fnW4vKZE5VpMM2dWvsYMOG5paR4vshNvjtaWVsC3
AFe9SFRQoc28DJjhdr7KRZYMLFMPL19BO5fhqdnSk65p20RUayUj6icsUCIH86Ig
QoKxYAiYoUJN7ZMSXK77ftiCwdjrf8t7zuzUUchFrT3lT8cLELigBr7LH5XWwJkW
O1tSp+QSeEqy59oXzIkewXuXiRy45OZ4DyVl+TJF9K71gvr1WpiynTTbGvR0VUNr
CQWmfZzupdATsY81ccp3O5DdZD7XL1TMy24h0ce2cDOYYtXRhdp5Pq68gK4fF6pe
hutnlRNcPOk5qNQedcCbeOgtBKNsgrVKnwCUImk4bgn8fXTJTgP4bHf9tfQxGQKS
J3Wk7eKolFi5flBsJWcbdIhVp3pLmu5TQsB0ubxdz90G6lCpj9/JEN1RzYsTi5wQ
52+UgapvGw3KYZcEIaKzohR+xebIEE+SAaeAka2KHCCOUs7EkeJC+0IOvnttOrlH
nlqU32tlTnkeN/01ulem3I3Wp2Szkc67/W/auHsudRZyp/3d4E0f5DzzBBqu+6V5
lAXk4CFUrj5ScJmB/ylamzDNlrvuFcciOVwzj024JFyJoSQakk1ctxY5D1dTnB6/
BPa33LhcGZgyRtC8Obu1SUjUj6pW8YtDNmFsuVRXQvO29iSJ8Koq4snpBQrY4aYY
8jfmGcvBdzQLgAtQyQ0wrXNj6j9P+v2eXx5PVYUmGsdTIvg1ZDhvvszkua8xDLMP
WgW73B4Wv2ZF8xTTz5WYjrxg5DdXTBGjMhp+PchXFY2cnKzaDS+A9ILGol4/VXaG
58A1CJUeGR7444h0gFyj5EgsMG7nfkqolxMEwxv6XjNZX9ZF2E5ZwX1FhvMmYPgG
PBVW5KF0HeTOBUSmNtZdVY03TOd5O07aZaWuMQYAM7i9v54TU8SCKyRecEZEkLgp
aOC02f6gwAQmTE/wMsJHAJd3hxILU5Y70KNcGMRTibNqbNT2ryfH10u55WbtBkqm
FIQ+XmnvjBINuSAaypqGH7V4FlIBK4Zq/a7k3zqxjl5o25rWtHRCH4tnV9+nm92C
XEe12K87aCdQIuybBQAalmrPsi048pLXoi6/aNGZ1GRoi9Sid9SAF+EqelIIxegh
JPX/8gdFwEPUi4BYy3LrnZjxuYzosa7QBDM5GD8S8oj8SgK7FR7IiPh6A3X4GIx+
7RBq44ad9ynL4TY+P5MDx8YSO0xpu2/UAvmYGqJ+TWAt4u1plOL6D5Lu/uWfhCHA
uc0amf7vA9GhEmL19kED49zv9+uxjOGUjtQdHfInSb9haZzds+jLBX5PPKWvRgve
BqqF8NnLyK/90AIjz60TqW0NlSFwuw5SsEhNoaaRZr2k4kI54lBHeJ9N70C+isH3
iVnasaNqFf5ExzMEWvcNqbTDMM2QSc9IQQh3GF24+UIHAPSnuTg5TAjjPG+Ji2qZ
iP6yTffudSGs4lVDi+eC3oJhHCaxCvhhK9ZGmCzPA0tOSkjY6+/JWaBk53N13SrX
w1Cs/SWa0GNjuhzo9mlUgOHJs+VhrJ0W+5D8U+jFZl5qbg9XZBtEAsN0fAuiBtgl
lS7aIVGlDF/hfn8WMEY/AARbC5r3dZYWGPVjRYFRzsDPzC4PBY6o2pit+/rJ7q+X
+81nkuFdJb/hqDO9P8GHFFEMc6+3y+50i7Xp79egchtMTM+s3cxAn2a2Jm5st7zj
ivhQaGznlDBHS4+Q72LEeJTptE5/5QXlvWJ+36mBj1MFyBFUzGawG0Yr4XRjZyQ2
D/zQtFfEkigHDsJ82zd4uGkCcUFypOKnFGBA7OAKgKrQN4VnB2sMZuKqRPzPf6Sk
00M0Kr19XdagfQ1P4Nr/vUCtvn0baKOvp1zbSlN7pKvOn7o6R/Mq0ULyuSIj3vA6
GrhMh81aaLhxyf+lyNwazL/tcqEhjGpJyXVAdJNYbZg7CE8sUuT8qNjaCEK77qs0
bux9c9VcfxSOW8hfxSsyrk1uyqfJN0290jumJzi2yLkypyCoCLiTbFuLDuMoNvav
PDfYS+FWR72e1mJdXI4UYHYl5QlBYHEVjou7a+tzoEAnsstyvhuSTwMzyBbKGx9X
pceO2Ag8YLjnam08vGMLIu1nFfkCa19PAfTXyf6ldb/gNRs3aTSUC4AbpsL4EwjK
K+uaNuCrUbCMJ4hVsYlstgGHWmFkvh0MbGgtc0pGoNvVDtWce+vjD8y5gR84NXCs
exAixsyxm4yr+7QGgx8OYaEBDCgV0zfINIgsC6WbzeDzQ6AGWfFGjAxDl7KNcfka
8++0eZ41/7b7lIzOaZhXxIXntJ5HC+0ftOawsHP1e33puG+MBcxXlHPDA7k0yOV4
ez3QuyDifuXCBN3aKmp3CQ80fbUpJFhkx1C0CsCGsPdlvmnB8ejlr2yl9lcYcg97
Hu3FfImJVaVdvwZID8oSkQkSYuDr6y0qKYyuog2kzqjaE2ZqKCeT6TzhEnHGNK3q
NkURfspjIoKFgfIFlG/qYtGHXhw3rvDX56PVtAEaHrZVg73ePxRQylyDet+w2hGg
Bm6fN3YDCNT+AHEbqowSu0mDZhbEZazigt4s3GQ3LM4uY6Qhfx6dhHp7LoPIauF1
1Xeg+8Qe58+/fm8pUFlTd2wBAo+Jw4JT67JZT1ngs3ojGCoSf7Arfh+Hojq2HRsZ
CrquXbFBg0QFgff69y859dzABIHDE4GnTTbgWDBiVXkgeRC7bSknTh3T+kfDUONs
g/wOYQlfbSWqgF63gUz7bGLfNRBCNKuPV7N42M/Plmqmlk9QKYrWi7pFto7t6k9p
6CRsCOxmPlDzCYmpsi3KQwaq/Sqd97c0w2gNl0FwqPBOBQjfZxkYdMczDrgyk39M
Shnzpf5YKGNjwxHWF9S6PMB9RHZjqCkU4MtwybjCO0uSsnoTXjSze+oLMH2VT8Pt
Fe9caC6FgupaNbj241gshcRlNIe7FLsO7im7QhRAje8VrkZYDfhdYg7/jrotcU38
U4/Nx598JFfcch7qrnhEhGEnpo/L6ZUgpb3eAeiUatkUhzWoBgK46DjIU4yfuF3H
eb50aJVLo13x3W5ixGrKj9ck4OoqoPGGDeooAOH8prVl3MRIZgWmL7MQ4Kz6g+K9
i/CBYd+Wax2nmvV7q0Jrb01HtCjK8ZwtOvZy4xi6Ac0W5ZmRK0t7uhrCbw0N3Ufd
1UclW+G4aSGaUxjF5uGy9+KgeMiYrTLYVrVUyb3iR/MvR8ZmMtwejp15MOR7ra7Y
D2BMfTV8kMkHgHALkHaNuU7OV45FX3BPgwJaoM8efEi+tD6+o1U9BiehrX9tLML+
t5v9pHLNR2NMMiZWtwt5J99J9KGZSHobbLoG0cyXnM22OCes0U5fHh+6Q3OY7HMV
YG1Y0LR2JktpYzopDt1AZEYVvO6dt7WTwofiT56vo531TCWKWSNsTCTImSpdrL8o
wCtdhLhuWQfreoNRf8UBixNZCG5OAxxFo10eizjSyG7TCh6Yvbc8Wae1Xownrsca
p7Eo/i+V7cMbHGGuSXmjbHXdn/4jvDg//v/8j8NiEgyVUJfkkQVIlaVYdNMjiXIB
yhcs1IMGCARl02Ui7k68IBKrbrWQtUI7lXedZ1gk7gDo6jFSyqCJBQ58MyRMHmL/
g/vudlpGs3a5xD8eAY8M2pHOVmxuqfIOKtUeouqgBoHESrkZQIPR94hlJ/z/7ZhW
er/HmIIjwmqe8AWM5fkABlXAc7DUbkEUOGpt/flrOQYuEBItsLWA5tAfouw8OP0o
wIgglTERWQQauVynEhAq1uvq7NzwIvIJLFP3gN/ple5nFoYIgLXpXqR0gC3ASmML
2GrwJkcvDVFSClLL9h9Q726kn8we13s0jWvH79v7ftKUwxv82DovJgRRVlcBy6lx
jb8Di9C3MDiT237zbdt+Hp+t7uj9vLAJvM2Pd9kgArPE4GDeV2GzWDHrjR0r7Zc7
b+jlioEIb7PRpwUoNXNO34+kk8dcI1yBdzJF5UcjJyiqR62VbBzyZ0s/OXKMhHmc
YaXucWO9iRyKO0XfSw2PPqzM0cCzotrsKc3imQOZVeNK4YhGpBHkiGX3PSGKU9My
cT1Aqf5Vs5dRlFKgZ8ExvbUftaAssmQ7P1xKvAPI3VSyVza7pJjVMuA43forBWpp
t1tJ+LLUy6jg784R9Eh552wUr74ArRFY1pxGH9SqLRJ9QeyEwObbGTg8vRnN+TZW
Qex2C9TPPdOPXuFyo9wPwdegapyt7IEwd0xfw2iYFXRHhQKwGREnFdaUO3li1E7c
vlOfQntXa9fCN9MezNC4fAVtmz9X9OQP922RtWZRa3kEkXK9esNV9HZeGQNr/dL/
L/tgm4TF/5Itg+5VCopp7f4BQGATHv6VDN4dxt8LaKS4Y3jhbBl//fMYnYx74WQE
k+dcRbzWkmZxdXTFH782zAmVOAy6Qc1TJ2mBccmkxesCGNkL5qYUTL/Ydsij0DD8
5kX8E2TefCoJD6EZwruOVIi8mUyqgV0MLOqDc6c12bk268xzgwsUpYg6Q+SWbZji
e7hA5JoHE7zXhpruWEE2GNO6rUFSE8E96TiJC5jmnvSrkF4w5JEkcAonSNnogwcD
3hOxoag/rRhrJ5BuuUZzE+9ldxC57hJG0oGbh82l/X96DO9EPt+c8cdnPA3wD6FA
pkPk/oPdYioRoqIiE52S/LBLQBQJtk4QYhpI0HCqXeBbKqpPNFJsWUSc95b0GKxh
Qx53bsVJmmlxIHFWZdeRa/piH0/Pr+ltSrLLJlQvbsaj9HcFO+8IvoY3jUKw6TzL
E06pqDhmYi/pUQFlE0UxbjD1+nd35HerlEqw9u6Rz08WqYZlLwSKA9sQI5+FoSy0
FgKjJGv0n7fmlbZRVq6t7764fVdq9+1C6r9mbE8kwMxEJCuQpUnBYFGcnWE7Wqe1
ORTLlwfu7q4FYSAMYM72uv1dLowp7DpX2hg6LMBKSMRaTXHXWIN+8r8fhWLkON2H
Ae5FjpT+eSRZfnMTYoDCicEtKnvbfbhkJteO/8J+cJu3YVm1VtDUa6P3PImdp3BW
8eVt65gwiQfYPmfFkUnRTcUXLNXYd3TZ/Vy6uQOeCSJxHSdX4CKP5wxiMrg7ASbb
REDfP3/AGjYlmGKVd1ASDwGjSaCB5Yg6zA2oYVP+wOz1K+F/xCwn+MTDh7VG1lvC
wW05jk4GzfwGHGmj/l3lkdif5cnhfODIbY1H7OcghgXJSk2fvGB1IYhRJfaJOz6A
bfmltHWouV3ao/X1DGj70QIjxsNo32IeTUqSj18bfhL76HNMyIt61AiQsnrly2Ie
Tt8ivgBiBV6gve4xtJY2pAQlNnNFWdoBPxh5qfAG3dKZYfEEr4cV9668P/1fPaLi
Dzrx0M7eSOy3wcvvwyErilVYZd3JpO/OfL5SE/HS+hHyQOwDUzjnXdjQ/JRanArF
t1ipeCnJZl9mk/HxFJBG3Ak41TG84tIxb32VuY82B3S1iBWBfYXAhFaRhBB/yuCu
A3JdyEk3nJ0vhtkdBEY+VxfWklilVWK4TWgqJ6CiuA0qNk+A9lIIB5rzY25sVGjZ
jAcIUZ7GR8KLEmGmI9oTWAHqM5asayVc9Su33mLfcgaJhNb5fMtVa2/xxz+RIFyN
NO0I0xn3Mewng2APw6hlmijryQOgpEgjIxNJkjdqLRIKfT7Guqa29v+prcrMQJ+X
BCTF29TgovUzqfC9VzAGqwOhR3sTy6lr3k/scDxVhNNsTXkc7KLEbp2den7CMQjE
yGHa7B49wg28wxV1RM21qnQLUjY/mkSUohnISd3triYhibdZtq3rPgUiGTyJM9sT
gYhJiNSf0cM86kVRHuI5Ebp85GcnaTArM18yDJOs9Ay7cg7HOQRLLW14P/Fkq9TT
6RycQRbuc88/eykhEydLD8zs7gcHVy/8oFfVARpf8QGE+1lZzF0ObTHvAY0f8A8O
Sf09gzXQa/NSZ8xUUAaFfvUYvUaRTefaYHqJPtUCskDt4mIWygH3NnP1Fvro2ItS
1L7DiLJZdcefV3l9lR+6wUpcA+EQSq2/OWLSLDM2Y8mmHUfPVk28MqdYSEziNRpa
kJnh8BnwIqzTCIkxtrsfckLcTAI1CU7gU4hJUBcu1FZSbyRh6tpYOqqQjOED6ih4
qn5b3/kMu8FSklS1b1tbjZYfgLd+N1U19gOeL1QH58k/AL9M0mXBBEsN7hSq+FUs
OVOgJIEikTKaH3tqJcu9j9yL6H1WRNui7f07KL8xq3V1upjMtCsLVRUFqBkbMjfr
CGHM8W27uT/7fv5r9QJdfWctZGnrM6YPbU2fJMLl7te85IH7T6TaPHAm69AfnklM
RUoXKA56VlpVQDGBh6TsuMVqBSocHQx9GOMUuHNvLisnQOvQnQSkn9je38GbJvpl
rYuwddn/hHTCaVbxPsh/HmDaCsm/SyckaoLtRrM7co0+IWwibF4Jl2qL4lB9n094
68/zSa+oAeiZ6HPadqVcyHGlaSYZZ5qeaGmP+dS3ux6xuyjNw2QlQpoG/WyySzQI
DS4a0J6KgpshFXLDlacenUY1UO8VsKtfybRc1WKCYGNQ9GoTNFdxhrUvTmv4rbmQ
XlDjfy3gidH/jUcnExyRARkTbGUAJMuIawDXUTsxvOwlf4Sk5mrno/Z5fShgqsi5
FYDQ2C5USIYxSwhu3wbmRvYWBR15tNR9CZz2ALzd9btfTuLSTjk1E730YTVT+hQI
CtHanlCrCWG0opJYgcuxR70ft8YHsQBwsF19j9sBqRt4I0hArcZQkfozE4KXTxUJ
eF5noBiM1HKXaz5Mnpa56f0pUy/KnJN3WP/BN4UgsXTGcVUZy7GbCDOWo2wTw0GZ
LTxn/y3S1Ks4PS1J2/w8qLLQ4dMhvr4I60FTp/c15RNz9gERs9xF9zNq/L1D7vB0
4wZ4bMw2tS9dBGzkoSTeeE6YvkI7aBteuPUbnKE3qKuJCJP39BZ29JtbGgMpJYsD
smZzHPGG2CDzw4Ut7Whij/gxlzVrJXO/TvNWQMYXPXvkjxxj94XI7p3cI/7od1q0
2ezjhaU/ymb5LaZLGjWsYgEnqOp1Nt7UgTGHiHNUpg+FblelFVpCbLf+uowBAp4/
pBgh0YfwHnhQCX7QLGoThHZH2Z522/vcJJ15/HquHF2f4zbkv2Jwq05Y+TJSJaLs
q3psdUb8vT469A5AV/H/UvyDUZxo2/jP5HNBWdpzoGkM63I3wSK6s/IE0Pih2tLn
DD5OTTwIBMuvKTREa7Oc5Ua5EzntgClKcQRxuV2/aAkg0U3tCL/nTZRU9KDsF2uZ
otjj+rNcK7TE/qcMJP/lOosuKrdJZOjTepUDo49PMW+rpq9NspX8eioTGF7SyP94
NE7h1PhB805go30SH4krsdOv2v7qPRIzkV+gC7OeFmesdoDFybW1h2I3PODlHZsq
8yb1j+j5py6dcV5yaZ9J0Chq4UYigPutnnbiiue958PXCRBrIcVJ9oFG8ErgOycp
LejKier4zhOSVmT+Es788n5Ce6SUxmhF3l10SawzQXi6AImndSonMmjNaWY4KMVG
b47Nt+9CKlmC470g0iNJ2QMuVBATsovR+8K7F3KSaws63eJ9L8vPwgyT0fjgViJd
BTsebqE6UTSCFVTFEaOPRYwzI+FUCxmiYTqgz/aCeJwoqucvuNL/Lpapyol0Q/JD
XVWtiGaDYXXwT8aaw3FLJ54tw1TCHthtIvegVm4tATTecICCDIcIhkMfwp3ViP/i
j90/jT38TSQCWkaq91btGnoZL59xPuB/0ITwA77BGXOtdSHJP3fsb2I1sW6X2dsG
EZFgtpLhFuYm05lte0LTU/ehaSiqbvuJNNv8+GliLAOSoYix0NviFGJBeMUp7bSQ
5SVjSRDKt5CDfdKy5Fdgr9LK2CoCR8fWRLEXkOjeUKiCuKedFsw4TQ8LNsZZT9kc
jNARkI9H6TlbHzISad0+yeuR3Iq6XlLpTC3OENmTgZ/aZpGuYWTOxv7p2fp05WEj
R0AiNOGlPQgD65zksmWQsofRMt28JgJe4iMd9djVuQy7TAw6eMFi7Jr6HNVbLUpt
WiSGeZ4XL21bFx8P2Xj0bKOiDyWpPJ8DMjkIU73PZo+yjX1WYeZoCbVE+D6vZbPf
6MNQsXoTfPt+3LRX0PJGs/7GEXkwd6vjiGSx1Bvf7596jl/RO7wf0CoBi/ZN7MfL
woOljq5F1Sx5EipMgNZDIumCINhsQVSv7cmlbAf3AovNsBqBuRqC6xoht1EAnOkU
d6+BL+111gg86O9/2dWezQBz83ZuzTAnOAe4T4KjQP78oECiZIHR3uZLAHSq+Ytc
HHm8c5CpXM6V2HcTEwVif795fGTx186Qv468A8V+jrfsqzd4RabZ4unM8zhloixS
Z6KmBZbF888xe3nD/riASKt5H/crFlqPc3G8xtAdewWFuGOQMnTLEphxnOu7wH12
3Qd1+FWKs5l2VHf6/uiPKib6ntMgMS/+3abjGwceJQ2Uh3oXnirDcpJnHBcPUOZh
j3CWMRayp9PQ8Khd83sp93wy6iVvf2BIUFbGoOvAfIYmPFlpLoBZNlG0tszyxWPO
NplzBceyEjtXv+WFaiXMf1X+mQivokuGd0YVTnOQbEGa9oOsyLEa7Fd8mjWAPzQ+
F//vkJldxuU6eTWJhd1qoMicRBcUHrhbLliyCWjbvQ7Cuv9LSL8XsLGy7XyTUt59
fhXXEOOtTvembqny+T8bk7n8S2tYNdOU6myk157/+c4o01fQlKifSfsmcqsw0siT
xbNNHOy7Bl2qU3rBznDkPIbCvnjBd1gzkv8jxTM+7eGVUe/s2wkOlscMMjDSaHR7
y5ZFYctrzcwyG+CUOf5thsc5+W8FFFwyvoMBotewbQFMhahCqacKZvPhDK6wr37P
t33Hc/O3Oqcs0M9T5TBWuj11w4JCbessAFjnq5hoApCQLVyI7tmUiSdYsCyHFJOo
t1bPpViBv3qPo1NtV70sEvFuwUtFYERQemZnb3XCrKQ1coH+r3m4lzvfU+XLbSDM
QAHZA1SP3YHeBY36bHLmoFo44nt3pxc0uzN9tSZEMrxPvEFdVNx01JVOh8ikUgp/
aAwwiTBZDh2AU2V5F6xemx+HGloXPKN1VKVommDV4ejwvDfjV13QJtqHf9PqAYlL
GE+/vRMgG9LYAjvRKpd0kEZO871ncq6T45GkxS0qp7R4QI7y/Qs1y2pU0FnsG44P
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ays5Scn1ZmCaOs0NyW/ox/Uaw9Ot7QSyg+2jzhhfrvSUtQ/QvHN9We4prCjpi3ua
qoBq2D+wAXt5Nk1hCKakvMrfMt9zA9uT+qYleQ1galmfeSrsHWid+VuENtXjG35S
DfMq33pT38XrXysRskVSUuKw4uysOeNXnDVR6U8HyWkjcicKrN6eGvwAgyE31Rre
WVgmD3Xe4Uyp3n5LUOzU1Vhvc5dCHzTDb+AJpmKiAI5E5MQdAULHjW8CACIG0+tA
pgShC0mti4TBvf5yXuG7pS3Vz2b3N71DQNFdOjQ6lqwoit5KJZig8ZFC6etm02S8
hTp1362Sn/+6E2+6v5cmMA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9856 )
`pragma protect data_block
aCHu67/QjvyL0al4V2XtnzivJ4yT8S5jRdhE96j0HGxbdw6XJ8+sSyeeB74q1Zwo
HEp9MbU4x/kEMFEP56aVv8yIraBZ3yJGBirClnpGRPzknPjweM4kwSJ/buHmbChg
8Jg8pNNyoQDnDGnayJO/mLFxq+Ig6v2mOxtERsrX+RzlBoqhVjmM09RD15r3EtKi
7Y/OgFe/i7ofnncVll2TjHbN8dR/GZbFnncty2uDcQxRQID+guR40IZO+NAOJgKL
3KgkwhpATmzJ64paqSFNiX5oZ6ue2cifMANlanXkbal1aLB8IwZOl+SOoz/i/k95
RhhmfO8yMvDTd1XutGWl1/pjEuvbkH+EuItd9oLHV9DETpEboWUGIicbC9QYFb4W
ekkYrguTKdkAhINuqvRImpmonU3/UPmlXson+Cdj0djHmt2GfZgfn3LvWVnDm5hd
fpaafG1uAlYtJ67j2tMh6WsMpogD/UgkhZ71JTJyrIjOK9DWOMx28BUUBLzdpuTC
ejLLXaFUB9UVORjEFH9TvFkDp+jqPZp7pvcMTeenZASd9cxoQKwSwzu6nxaVUMAF
2vZ+b4TDQsrztydq0GPMv+OYHYXdsKm/YYUKQK57u5bQxrGGvyliRBNBdTHm52UW
uibAnmc8kYtPRLz/5ouYS/1r4WEY9dQHN4UesyUlXKSS1o6KKVZmHV7BP0EwR2Mu
xxuqXFR+6VzUzQOSYOut3MSVn7hPv6vN2qftv6f96D2UlT0n3AzDBIXsucfR2ss6
ifSi7P3G+SG8Z2GjGrQKk6yfbWztGm5LxlYlnAJuuxzLQLt98lSfANJFtcC/KdEy
8wCPcS2zATFlDZHNPc+h+X94XXAgOKb6zp7guFevLlvtImKrMo/Fk/3AHeoRhOpp
IRxrK5BfgBVBH9PvtQyeCEwhGrTO3kSyoyMxYTsYIEjQYlXRjKGlnKtMcB8RUXgw
iYk9nP3JevRN3B0zPF74o2oRs56t6oXhlEqpFCFT+VTA+xHMaXyNsLA4gFfGZdjS
sVEAojxFS4gG+PtvA/wuFEIG0C3r4NjS/eaXG/poP0ltD4Jv4E5I/rQwcdWusdPV
hbewmLVXdF0jT+xhO88+2pVLCwsirj8RQOzH44+eHweYAiBu0cTToWLoyNJLPYud
/AZXVZFvv8VCFDeUZxPg3/8e8UTNjL/1P/cUlLWvVPU+WssE4npRunOIICLV84h+
RvU8nfTVid158a4Hb4MHXDzkM8RPNUC5hScPq1/F3zXVCAwNIaYXs99ok7gRuYI8
atOt1HiutYWWtfxRFW+Xbo9u+Mwd/y9V0y2wT8P12s01D/iiEo8tI2lQVCvUfrUG
sJ26y4P8d78BQVq2ByQcK9OZO4xGj4o4955YOesz49ca4iRwy9VLiF61FfPFnmyr
Wz060fodGVPE9xcYxtT1Ap4aW0OTOwbhUd/pPGInfENFAnrng4+O11Lyd5Q/CC0c
g4LZXkrFuuHs+Zn/7nkkMJU66LAPgTAubmE3usA6Otsoy9MYGI4ORujR4fiHyMsK
ysHdD+x4d/+EywVn1icU9lRqM5gPw5CtQX84FcJZxPpTsMDSHe2hyrkwPL7byUzi
K2j9IsehTheOHX9ITlOLKECYdszk4vrqUq8IsvPJQl6QlQ3Lu9IZ2QjyC0E8zP8Q
C0JI1C7VrZ/xTfWAySRyFNxBG5VR7IEuwLDiG6i5GV6dpju77QNsxs6kcA89jQ6L
Bv+EvovBX6md+CSsmvKL0yT3rIFAMgNqK0dr1NKdKO4zMc1ApLvDLvuiyvn8Y+gh
Ry4L7AfYya1xHu8Y9cLJT0hYnYgRCGsbF2tOpxUc49t7ZHkG310uikuvI8zoUQgY
KIB1x/H0IvTng9t3K33kFqpzJvRbemWPZsu5BsTArPqmEw5kISa6Wi08ZNjGWlWv
fR3BuVvCFxcgxJht8b4GkiqL44rYm0qayf2P6P7Bk3vCSvMaKilftD+dxJgPXNxe
7ysf4xWYWnncp5etXAUG0bCv4gmyowBhpUCXcDIOlEpdMfltd9Sc094ULnbtJE17
FjxAquoi3p+RP8E4TAgmbj7zPTgr7L/SxAQlK8aJQ8AKDSzD/KOSBYsJTsuYZKUa
yCIOQqAvgOGVdjmP79ZoIVautwKNOlUWAleFs2Lk+05MQpL1I6LKXZuqSaai3fKt
gqVDq52Ql/Q25cvPXnanWi/OXKSSDPxrpSRRoKtDimuF5RBdhAU07Ny0Y/k1uJ2N
ejWAzhr2HQXomd8VoOlk5+NubDcLZE2iajJeNH5eVHoARCKTFe+txkbKPnU8FKPD
z9W1bnX1HVsPvq/JjunrBO3YxRZxZY3EFOW9nY4CnpMhE54e2qv1wvj+8yQ39Ti7
LypOOaKdLUeviIWLpEHb+KWY7uBn/P7D0E4Rp/tRw7zavn8YjDe24BrjuShR0MZQ
xnGMpSgcXSmVxyMdZBgaifJE3o+BT8QjczgcLc80SGF5uaaLU4dT35HMMVAyPWnO
dijVt2m5xgitiKUEyPZD1GVjjiYm/zFZevFD2PzKzIaM8cf8aZYLbS4LtS5gClEH
crNrl/+6NbzqtdKyKi5Ch6CnyLUkfVHFf7fWvTa15jDDIPo0jvEsV98fY1pENHJV
7AzMPGNbAnXVIdQSaiixT/NIgArvvGin65olplm/C/WUyPk/mxqVImRGE0BfThoC
yy+h93vJO9k7E4YuJjGtsA6vy4Jj69nk5fLgm0NcSERsL4ANxN1b5kvjIDNeFVdr
WrXqtwx1NCN/LKIoTcAIgRdBZ6mtzwDDb0HO5WGSfQurL9xbpRC+JNlsm8Si6Lho
MTCfDedoYIc8P7K92AEYhTVjevbbEAam6DbQWtDoMbnqC8/gtcxIfO2QO5pngq7/
lcCLlxcrm/qb9aDFo3OOo1c3PuCoa5OBem29fPgYICqCugJofQ4fLKGzJEwIlaff
p1QrhC9ia3CmIFajjyxIAEtp33T6vWVfH85NN8GAjR38aODsowurbsSsQxv5hQbg
QKacyqm98lIAXnFI2NnGlewmgTHeo2mxCwbeCTqOkZw1e1rsSTZymQPeb73QUn6i
qnougBnjyDW5I8sAFa4PoHTP3bPyiGimyZUYJcKx2cU/dHLZm+quvuJrh2XxAreO
3dS+9FsHmvtIv2HdVetVlc+rNFJ45lITpsRG3c0ySbXZC1RfK56mEpbhC0sWVojv
DwAimWiYrJUIcPRRidBswZvK+iNHSA2Wu9i0Lrzvq5miMsMCOKCm3djJurOaMG4T
4yl3RaOchKqaDuwz8tZpRQAacr4Nyy5w/8e9boduD+J0ak7nC1LyT3xVGnnABFfm
wdA/zUIE8eMcquaDhlVULl7uteFWsk1xZco0+4tfMk3dzwUNY15Op32p9EBsRF34
CBHFvUw6tAs7iJq5Whn0uvQaRqo5slA8ZLD/POMMKiM8ZWUf5ggjdht220wSBmSB
IhfOfiUC8ej8O7a5CeogYJy5Wo9vzODNZvTuz6L8WSCX65se0RZEZfxIzKuwJkq7
O7hda7EUVOUzQqONejsKxMttuv0eHRXtb8Vpf913vAOWgLLfnq8N+GU/+HIAaHjR
niShyHAMBb8eyEdWKHmJrDN36u9olvJwXMqC9RYHbFd7KJtEweZuNlUWczMkTDHd
MDu3tWqdfRnOjK3Oljd+CYaeMgg7zDRoa95xs/0h1zisuihVJRhQMKExWuMrUUxh
ssAhaCaJADIPjLNr/Gd+m8dYJhmd+eH7+VVdBV7Hx9yXwoiWanrs4C+7RSENtSUn
Ze0b+jkodfOlzqj3j15vz/RPQZWInMPfNpXjGfvIGdVet0aIw/fuq7ON5cTdPqty
l7d/TKmSZFL0nc2BZ9krWa2tO5o/t/5voFA0/tdEQ0a2HqIq5dFcMoxnD9jdrl0r
jkUqsgqZlyD1Xdmq3fgB9CJiDm1UWxaoYh5L5oP93CLxWD7Zs6bWKj0dCWD/XvX0
LdvRJL7ONMCo4lweiyoAqumxrMkeH7uln31k188hKAD8A6FOgqHePX8bh7T8yayK
u7GSM9JYN8a1QjqnOcWAOxPpNk/FagLEEzPsPtD6YkpwETgNjIV74xdeUmmw48OV
Qw93JvDmE13OhITMSwc/i3o6lthBpGZGywpEcQE4M4G6DOTpAvMrcuvl+5cpqtOt
Xo5D9N6ALtBzuHP0OjpKgljEWrlbNcuzmc1oL0qDJd7zMSWFpvMwuOCw68wyYcaS
FKVYs9/rkh77nx+NyS9JEAHrMImt/RJxdmxS32Ju/5N33CDsBGuxOKlkeHMthNg7
c+6g5S+QaWTjr+DZymIrRYQu1USWx9oSG8EPc5+ySOGPwXP58BVBEKZ3KLs7VnZh
aQqodiAY9PzbqvMkw9jdNcmEE1hmKkMMCuf1MEFNWw7gPKfFdtmlnHROGrP2dWfI
sJoFrlH4j3nLJg+8KgUxWbQpb1HDJY+a42Ta4tuXsdrYjM7wumCkoC9JiUNx1mMp
2woKhZmgwS8CIBxbpKxHp8bdQS4k4v4YT2FgQCaQWIwrXLDb2i7/YLegk+x11j2f
CTRn920utsIopTTrdvExgYgtn0Q8s1tR7/ZsILqKItTz6nZMFRcA7k5Pf2gh9L0U
61LVZMwrMK5gUymOQ8vowwDfUn/fMHlyApLDKkejosJBHFbrN2capDjTzEZYoqp6
+TRTRWxf1yNtVE/O4+awd4kIRn4a86t0vU+QtTVC1XQQ8w8XZPsJnf2MBPYu3s4s
/qmjT4SJClFY31I5CaY5s+jw4/FERP6pSbFR8KVvN4GZN2Oyw0VNPofwSKtwlOM7
TZtMnX9uJqXVb7WwhEMV6d6rz6S5bNC8/xTASjrdLPJ54RWXeNaZcSCi2VdSD9ZZ
dJiRR6isrfJ+bpbK7yMln2ppIdIOAosyhzjM2YP3VZZy0vKyWQfjnUa+5/qPBxHd
i1t5niKRF7any3H096z/lqhMR9BAC3bE5zoMFcXkS6DK7c6AgTmKUtBAzmz1mu5D
yg+YIFuEOCIq6fteV2Fzttg8AXim0cE2SF7bQZIBFJXmY/XQ3j1d1qF60cnadLAw
m6MzIrvAM9sFhZty2nvR9eJe57jPuIlhimQE3+e2ZE9dDTVvBgBCgvGCAzQ6kWs2
+GPRjZSqGsNeH7WUNB/VbL09t1ODOvEA+0hl5jThxwG5DvjQxf3Y8vMDc9r6TRr3
YtufGVrRRg+vNrjfFGwNg88b+ZOKphfaS7z2mqTYJV9OlZubhKVCAdjOP00qdb75
4W+J2V37kylcMThk2KUwouHXrKVfDaBvi3cFq8MnKIYTW8TPRSG6S6YIOLGbFund
j/Ly/hn4n6Oq5ogMv2ooDpw9oaC7BCrrmXuCPQz4UD13U4U6l78vEKeJdQgSV6oW
U2CFDve3wLPDyA9fqpT0pPN7Cn9COLuJP0+W/6h5YHDfJleb9+y6ItIpXhXa63Zo
RsmP4n8K/69jwhVCbkshlGhT88JyvwOQzV7xBQYdQrI+oD0/cBmLLxAzkGTgs+Xq
Ora/5/HS9I7fC/THiHvAXcB8X1/S2mJiQRc3JbnthVrNyprrQpya54nQtItSeKdN
yF7OhdBUzoQqhrVKszhwL3nL6E8nI8QTSpDBHn8ib9C758pQLTevb0TdyO92/egZ
8+oXfV0csw7AgOPAMf0q0p2W1irjNbLsKUxv5LBRkX84fdHmRTq6yfFEcjua7XCi
lPB+F4ER/W/IQyMFP00yCZgYScT0AO6pXTYF7qQ1N4PGhGWEp6itN2UEFSqHtUBa
HKDD2SQRem4HuqYjrqY9HeRO/vTRROG2r9SHmleEzFY8lKeSepXJPvpTdItAvRNn
9OfrG/o2/OgT78t2aAsSwxigrdiXNIJ2imMWsh+MQGxvF4YZKDyguihSMCXMghDN
Y8j38CjnJl6u/JRXLBTOEwfKtCqruhKxFvSKkLjNwOdY/LBOWsmtqFUXKOj8rcca
DSfmSvGimD8oV//3J8gVuFF6ScgKiB0FJDaQjPHWnu7xCoAKxWzOzn9EPE36E6dy
EKeoOAId327CcBSkgghYpPtpxkw9isIHzaamMXPmX49/3vNio/3R1I8IIKZaoT+L
rLua7m3xJXDe5EsJj0I3wGaTW7grXfQ5+RiExiYll0C61IfSvb3IPefvle1gLrBA
bLLX9RKaY0K8Mw4/CPAFvdS0Bkg4lukpQoRYBa51G5k94004fhx6DoxWL0me2v5j
ZEq3VXUZglOlJqgF4juWjelRVw9dTWLfEmSEbdP/tuAswJSPi/iPETWmziHBLlUB
Alo66vWburb3/rluCBdftHlKpnyf9B4BzCBhwHskLq+EqBiFpcaEM+ogEAMIt+3k
PVDc5jM73c4uzh833h3GHEnNBTmcszpd2rEQwze5BGijKJGLQmvkWZpPTDK3a9BZ
ydwt6fK3P+rQXwMigXm4VbOF585UJxAo7s5RdI66V9gL/FCFF05N/wpx3/nNXd5h
bWs9vcfOUPWMahdRl0EtkuFcqSmpkRNRodCmNnzoqwGtaY0tE8KkeNBf+z8uvu9B
ezdNCbMy9uSmLkxHQqK4jPM6ouqU1Dq9fJihkwoPdppdjPWGrGpzhfZLlfla0kif
8PCTjxnbp0itkynMYO4DtpvuLlQWHMYX1DtoO+tjU+GeKdt+iAwQgnBIAtRpLOXO
flVnfq2TX56aDLytV06j325lDHEbzlwz/aJOBCUJhgBqtY74uEveMmZ8t6y3vBeQ
gH7jHbjEe6A9NoboDi5RX/QljLexYKnXqiO3ZZmSy++TbwB8rhYKk8pZ61aFd0PD
9F0iXTO20omF5cS+36QzYu58I/yfZU6TjW0FCmM6K0gr2dzfX672hnz1NpGcibH5
oaWBQjcJxZhZQV1RneRcBVPA0+hvnhLceyMfyuIdawov3aZQUhiIhMTLgoqMGwSz
9U96rjYS9b/PtyC/Dv38Ho+LF0+6Q4Te+/vVH5gAjTmm8tEIsXtpj1/6Ge25mtZx
hsGRv9J9GP1AcSQM9LRBhFoKhKddRm3WRKMv7Zr1E/B2U9otdsd+SGtlCdKAUSYy
pGZYSHbKUR33V5kngeDgz16/Pw+rm4sxrtxVh9DgiEw+fBPNRBIbwzQEvrieM7RP
zUyYwHxxi1CgHx9UyAsm1WWsZyKVRESDDi4fmRpdv9Hk7sRSZs3trlwkuzcMCOIp
leGR6zQqTgEupbNGDQ4WHpe4nKMBb8G3ANFgXSp0rZsZdxqXHWFqPUm28h+eJKEF
dRjsc1a1J5ZR1sjsvTWbBuGjIN2zk2Naodd8y94M/eeEIjv4hK4CntUqcs7wPdvW
nrVhftYotbkAWuT6wY5m7VrBuPs90GKRKR62NSobr1LujSSuR1ApRKkWWnsL1+oa
GC6MDSoSI85jPbSs9ES6j0hXvU08Nc+rFar3/xDaGlgu29yCVfpl2+DAUZTWW+8w
FOp4scouE4YyolDBx1bLaQKjTobxyiOZhd6dT6gazWWSgBaBk0RRPekNXSMhZVsA
NKSDbRs9YioMkwFZU6+W+ruuU69MCwtN4EllwHVnMS+Hlh/4Mrjvvg5TtlLNOQcs
qI/1xzHGYPKsMVF13Tc21CYeac6Zv8Xir/3ndQcMYAehAnHIAK4hasLeDSEwy+7D
60X+LYAt5eTo2KNqkWKJ1HTCeY3AteK34VKNkN5c22VMj737JCDNfb3x3xXXsxTW
zH+wYJ0PHiqlQW2o3yTM+8zkJro8xveZw5XSSrgN9YGFas6wsdez9fE/LSjDn/ri
oZ3MjQkHbDeGPWxXNFaibQywpbC6cAdFdzpgPQQh0di5D6R9iqxhPZnyQhCE1SYI
ZZ7PiZ3irGWEan/IXhTeuy8mKwVuN44LJmPWi1R38l6NMlrqrHvUwY7VUbBzTuDZ
3ZtcmH8XG7SLFqW8GYTGlMpz0jjYrDvMAKLsGXF3j867mHZUWf31/oiEt+4fk5XG
ClKe19y7iPSnfNaq2TdTyF7UMX/RYSe+0MOqgt3VTu10mDVtoX8l+fOvmnwsSU5o
OSgaeu6CiVt95edlda6+IrTnEhYK046q9O5h+0Rnt7XdcYGfUfvx+EgE5bnI305c
e9UI79EPYauuBmkC+v1DoF1YnjoWXQhjGav95WKNdtPwmz6FKdFNJkhfmxGQgkbr
PVtX5B6xtFL4ukTSdLfzWDToPoKZ/6bTf4AlEc1uHEPcJBi5OICyeuzAyflhK0R5
aWZttGg6AQ3/3cON0fQ/X8uJRqcRbmTwEAHLIbq9CSJciBXQTk8ew1FNOqmFlMQR
ABvPVZhA2qVppB1r2eHcFCqx5yq7xw0nfXk1cNLQwkgRlLzewZM5FH/pRliIicVA
gpxSgwwkJSYbwC4yxuhU7cxYfdKJ1Cz2dt0s6BG340eClV5+fZ27NG3yKqU1jZPQ
OVx+AhBFQm6SP5CbzB+JNlI7ylr1S39PEf/pM+NKfaE2K1ZHzZJ60P5znnast/tC
NhJwocg9du4Lg9uBYPWWVxcIs5ihZYsfSA1L6iVFvMVUeKCNZLslzILsiqMltEOx
25KXTADlue8lvxS9tPX9J0wSZvHaYyDAk332VbPh6MTzISJE9Ps1DM+ul4rewv7x
3E9+cdq6AhdrHc7jQ03fvvrqmyAzJ+CCiUTsH193yuaNKgFn+RFy8elSDTN3d+x8
i5csK68LCQGYzFFh4+fQVC40iYOBDODyQ0onM5DKm63HpGrudPTKLO6vzorhrPae
XUubPtBdGAcZf5swQYnhYBg1qDqfz8ufG6RxhTMVP9xO/B7xkqLFujK/D+KXjaUp
sn+MDtRRq26PqWWK6TrDkhXXg7mEPsIFOJOtBsceP3BZuP5WvmZDJCJXoFGF2/Pp
o2KYMDp4Z/cDAQSFE954oMB+IFTmm0lxlpK4u9rdWzbwLnnLfszx7wp5/nFQzd00
Yvy9vDu1L9+X8cjvxSB3UwtKEYoSFo+N3OyKyJOOHRvy9qZ0F+IwVPS5DQYQ5mvD
6/MOgMpcvoXYcONAir//H0rpdbvhsPYbVCaXUJa53n33rpFxgU3YiQYWguxKwFHr
JSg0zMV1M3v4Afmr4dg6BlShqAMGTxZgjnVeOvlVe0U5EM0pAon+pL8lVznSMw9O
I5qMGPl0vfOft2QAUbRyHPJ3J0x4hzLhZLA23l8GEZl0b/pFJGpljo6Oja5G1pcg
X/CusvPCF9GCG0v67g7tSu00KBPCVaBGaPSVdDaBUvU1Ve/TWErRhTtvzKm26FSu
fvAzVhE3P3IUBadOoAqBZ1HI5Ced6sDhm716RJQ3iTIN1lHi42BM992OG1NjL7Lb
i7cddw67sSFceF6VmbbfNFbbAaB7G2GLk7HuZOCNFOJbT+uttjwMGaIPIOCJOruv
zZc3i2A6ZKkkJkzIjIB7y0rk3Yl8Tbj3jQQy9zIGAB4v71Ck5goOfN5Ws0uN6rVX
9AIGKxcVHVgLUNZ1C0M+NKjj2LafPVN4kDIxAt1WL+N3VDYcgIp/glGsr63W8ewB
xUvQbt//2bDYUQUBMyf1C+uNjSfMiLGtCt0eYLKxoIz6mvcZQs/2tjeIAmJnXsYG
WtX+eHD8B7j5ZiaqA/5bI7lD+vCjYZYHh5QfzHiCpeJ39s2iK/Jd8YUg78ZqnYCb
azttLr943Ul0ROvkpb4LUJ9PeHDEoL/Sx7tnN6CKFuIPbkFw/hkjphdQTjEtfOtg
L6bhJNjQBS6AqKC/nvT62Ax+njwfvA2kHn3u/ZJwdpUnhrhTDEyQaOD2m46Padba
rvvqX+ik67IJ65T+w2iTDu+EPi18TNLgQ2Qy08Q0GurAsh7/ElXyl0d2Ix20N8sX
uFCUJ5toAPw+TYME7m6tnVoVDL2YLTwsgqNWFLZyjmWxujRQN3JWRZrGtssn5iH2
khqXi1NjutrCuauBflkXyfsCgQrqDqMY559it9zPBgDZW93FEAEFrCTOBi2UMlPN
eoN9du4Jx7UidqavUFMG42AWbsN0qFR6PxqNWFQr5xKLWtKDoInzD+x3UlH4MkL8
GoZdz696a4aWlHzWfcCndjfD0FScUI7O+NsUxIqU6lQuJM49yf1yVkzt0NnSWsfC
yQinQ4asYaB7DzNpq0m8H44ITbgld3nIRDM7aqwX1CBeiQZxCGZO10qUaUdoReuU
6Xtoz82DhYTzVQXBcjZqGAEc1CW6nAm5HrjenRl+0rTfEFWFuGOoo4380fDN7mDB
M4SsVkFbKrqIWTIC9uRJnV+kILA7uW/rmOKkWTPUrOhSX+feT8NxDFROkRUZn1td
px3OFiuDFpXLRyEefG7Ci2mbiu4VKYGsJZUPDvrmNKHlHPzhAhuyabrKKH83DF9C
b4JrulZLYYJ2sf5Pj6ma1ZnkpyOwhOouMraQuOZUKnpE1MWzq2PCKtFq2x4Fybbh
lqyJv6Hrk2tUD3fXyR05ncILrQeOfWOWbEt1NYMKu5bDrjOfIOKCv+GaKgHhlKyP
+gONWlGVFqbc23hEkzWHQw+C+eUD5P2sXBT+VReq7ghH5EtwYcFLQ5ZsIsvKDrxF
baGQXTKo+6DPEXs/xiCydbH2eblf0Pxt3Z3z4OaghaEp7+IeHX+yefLyTrkDnB50
DQH8kwwBCcu/IHvLU0gmpDXzc+0kwdYaTySxYLIYPccx+NiIA88UWsQHRkwMXbKB
DhU8msGhHE+wMRgPxLiWswoi/QLEos+hGj4ltYqBjQusvUhG0Vey4f6YXIwGPki8
KCm+HpBHxYpf05QiE3EoG/RCfVYL4I5u4wR1sji3X5wkWSlAbeqSeKdMmYYGAWXo
bQUrsUgLsK3YxeuJ1tREXGhMV13wrlom0/2grh34g4PiN/S9yzcsXLemJ7G+aEV9
djjuK01pmbHfLm0TTiw2JL50TO4UN8XkSD6lX1R5FmRl1eTrFh0i8bPmUwgpk9V3
QeZtE2jous7NPJgXglR5/M5SpTcn6JvoadmgTX4qXftSsEi3samZ8RWOQNuQuXIf
QLUFVfo/pj/utcfVNDw+S4xIWWMgeJK65AtS6XEb0e/3h0vCQ6Y/AvVVP5USAczt
VwXKQqHPHCysm8xlrPotsP6nqEgpKf9f/KPFtB7ux80X/Z5KbRVT8Xyr/P9GXHza
+UjU/LGQOPJRdDRo/catBNqRwwPzD2vtuVvCPU6Y05KejCt4l8FuYjbuoRPffGbq
rv68OVGYl6r8kJWx0LXzQuei+BI5o2L5BYE76vdqvlDV0xhl6zzu4suTdLv6PRzl
0m2LPatmg/q5xQryPTmOVbSpIwI2i/zXezf1MvAdfaeD4mRSMoVCL9geBjwbYk2t
ygEBF8Mq2yg61gLIixDvqd36UUUQ0qNhLbQODc4IixQs7QSHvcpmk01IKdvsrC1V
6EDl31APTrm5Cvv/t7XoowzcBpNPTeDejZM+hsHPvHymZSonI4Gw59/fv2BB1XHT
2X9N3GVZOnUdZTsihvzH+TKW6z+yA1UXMdwGGkG/WZpJj+98JX1y4Ujxiy0lRhrd
2dUbaYra0P3lIt2/1JlqelY9hU2g9lrH0FKQDN6RPnNfaMWsaFHjGjGolOLFk2e6
HHuZM41NTO/027VKn3WnueoBdkpD1stSPxezInqyI2wLnDTChuCPx6GOu13gzpX2
xgde1qN76VsDBFxyVQ6xjna+4RhzLyPWQzDX9XQk9NKaqsfWuZ5LAz6oeFZlQENp
KX6bFlnkay5MnCdqo6xR9zj/mnI8DJ0bLpOrWNNe3itzM1HsWFHuFpzQ5Cskz5bZ
HgtdH3CpH5+iRNLMISQPlKBMR8KfWFbws0g4v+Kgwptuoj8gLyThhpBTQauaqnaj
ptW9Smky3Fgy9F0npU1PtrfqiJzApo2yIZbFijr7GJRGMi8nrQrYtpW1+Wyt/P5j
aPLTeRdvKqtQNMHdHh9pVzf+tPwECPP1XbdKQWUeonXMHJf6hDu7C67Vb9ux51JP
wnE58d1NNF6oh8tgt2EjU5uDqv0M8Nwak88SbGAoKgNWkCi6MhV4Ag54e7WTPqLj
KGaGOShkjdVQSCcGuoVGdou6ACzGHYF5VMGURy/K0NEIQ9ceZVY1GraNed+iP/yZ
6RY7XdsHXcMwIpq3z8PVwKNWOWYGgTlzaZiAtYVunKTgA0ANIMEk5xeJcxxwgO6c
u4EHhNEpRNn7Z9xM+J8bTzZJmcIeoyv0L44ug11/7lBfPBwlZ3sBXt/Gz8Me3oB+
Mlp4VDPMPx6o+oM0D67h2xprYHsR0v0DvcDfLHg/nHflML/iccsvwPrj2mDxpENi
Fy/6NssdXQlP2G1eyqOuYHJWuTtvGbHYPKyE9GsN8+QDz3Iqh5z25HBHUa9sTgWx
8uYAMO2Ft4ydq5z3uWfJtlmVX730Be49RgLAbR16mk/qetiLcYuMQOfd3C8EAy0B
Pwdbw9UaRm7RsdE3BkMQ3DxK3aYEdw7ZlN+m/8X44hbBh6mGkcBH0QHo4onQwKmQ
1yYLuOvoCWUUzL/1D57aU7Ymky5mMA4s9l1gA4wJL/1pAGjkS1ttdmBaD31cORMB
1m6XiuGt57ftJZspFutS+4ibzgVo+2/kSAPleGgOZmFL/y5P62vcNuf5oX+s1UNX
kIwoOY4WPYHBrCsVsRQGWpouFDczhG0cHNz5V778Gyc6c2ftq2aguqfWlRhiJy7U
f5zMulyqhnXiW8nQMZhgw9rH4zE8SO0yjwOR7IFFjj3OijuHSKplb49FLCWC3Cr9
n7XS8eB0uzh533KVzy365hgZt+HYlXZMyraXZ79wewshEaJkH8BNF7ViJtl9Hb+2
yyYhM03JY3mlP/kM/zkqC7n87PheQ2bUTsA+uOdIVPqUN9ZvPjb7pEp1W0YHKirO
XM6qQaOgz0i7DInQAWJIYva7Cd2Hifx+rsKGX2z45tOXoRDWjZSbi4XdbTs6IIgf
OZGtADOE5cKcM/icHbXjB+29TGcGjT72xHtzzYHdg6tNHbnqPSyIqY7vzsK/JV7g
eS1xPRq3po47VNjw81ZwAOnYl3VDxqj/ZXdXPUVCeb/ro2c7VDGlRN7EG0ml23Z1
XmNWtWUF1JyDPC6qol0fuVoVv/H0qb0682HGK0FOKFOyaMQcDjmg0XFJLVU2Or4R
UwEAiE9QBsMlnLFPRHhmfn09B8Xr92+jb527ktFBNrmTcy4utAq61+HOG/NXXSlo
szX9ndwlfd3KnUapTqqPbQ==
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WTQetkw7vbLYL65uLIbux7Mii39m8BywXh4dsd0A7obH6UgbUBea7es3GHzJqIye
+7/lDbqtkhJVlnk8IZJAxIu35HCWAHV4fieVYGQkUunZPNfinapdl04mKbK8MWOf
zaxIW7yUrXMHn0ZdndnN6DvVp3ajLn49vgQanOiuEHuOpG+lGSOGJBqW0d4Wtsyu
foHkYz/mQJJNIjHMKBIMgIWy/HJKpN9rq2bJX5CXsTwQaHb2WmdIgJpykjlAv4Q9
vKaBGYpENPNQkNsnsOShtj7H5ip64otdv+zFTn0Ku1c+JEVPk57wPSDlxAGbT701
ipjB6hfHJZ3SZZ3LDjWBoQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 656 )
`pragma protect data_block
NUJXUYlzYDjRmIhuMqI+tygFGwV9DnEqYbtCUDkswPEj/v9rGG+0SX86DWv4etsy
w0ckS9IcGAc+WLZVAJsGddNbd/X4sZt6rNWG6Z+ceeZIEz6JxfHq4jWhamOu4ybL
NiiKYD8djqn5Aea55dl/sXdXVVEmOh82TzpKj1KREBazrKdoocRLJ7BQPmaF7ewF
MsFol8ZYg2inKnP0oba0akeKMncHNR8Iuby+wyt/evgrVjYH9ZAp+tbFN8tNhMlX
t42XaxmYUL+yKAdX014XTm3gXV/T+Y6w22TEiIj3+9d5QL6wDn/6VrwXZ9SMtXJK
sr5FGYT57eJnpmlu7VFSnVfv8vspjH6W1qxKMJN62ORicgY67SrxIkrzhrXg1xbn
QMT8F2qGlH4Tx+Kq8JDANqurcrILHmGdPQXIyRQSfgbd8JQjdA56uFJv6uaMYyIz
cYoje+kRJWwSP69qrsoE6A7kS2WIE90ieyL5eOORqgG0jZ6h6b2wZtmcomFc5oUF
B52JxV0ztB9voqx8uLGvXX5Kl3e129U3Ea3yWWOYi0a7mpP8INBxZn+z0U8HBsQd
E4sxG793ah/GwU1Mlg/CaBBqFeyCW20+8ic1IWaFBTxM3L/ZolzhI3u/dqjh2UiQ
hTv/e98FKbkb0XLLKLTCCBLuaDfKgk7vahgA2TGK+rzoSDgu+5efbO6ngy0ibE9G
gDwx3RnJF5hflnUZ4Wsgmpb33GIpG/ypz4hSYHkvtPluNR7Ihb5wVBYKycOuF/oB
C+vP1y37jd8JWpVs9TO4J+HGuRTvM0n0ltjNm0jZPu4v8RDH5YXYfdkMrDuQ47b1
Z7uZAo9T2ICfDHO+oSsaDoHsB6XPqeiOHwboNznppWc=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lY0yOVMh1jTNYOISCDWJAUmW0Yul1Pl7pw+jgbfep3Dm+kg4Xpo8IRDECI5FsUwe
9Cgj3inm/fsG9KbScfAJzT3EWkfdXRFTHagk0J6zi5RyFKrqq6rgyKAmhZIxKRAR
e0PRew2jdopW6GYZk1GWYsfc3t+TLWkhN22hzk92l5bKuEc8No5j2BByDL4X3x6R
K7rAC9+71Tul59BB/D9JBMJCMaV0zTvnSQy4JqFUaB42W1bXzVsA5klEUSJj26DZ
vaxwTkBTmrKdpIvE3go3AnIcN/8tMEUC0dGlCwXg77lhHtAjRMcVTxVGGi2plQAl
AI6UOlgzROiy/iwtwUVt0g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 13232 )
`pragma protect data_block
MECq7EDHQQnpb/aRa2Y33JQN6xcnFGb5u2llydoCzz5RG1X2rhyylm+1U+aNNeJL
jkIb628XnFAMApjx2NgC+1RDPprjlut6RapVlEzTZTZRsuCPSXAC2QU5yR3LjEnx
zOtP8naIwpyG8Ca8RHCUj9T6Fj1/CkxeyF3WnVmAm/DLDPmuKzJJdRu8kydTvuyg
hXYkFj35wJQoKm0Q1dVALW/f+MQjkYCLH2cqNZdXRSIMupdqomkiMAgahs8MAqc6
av1gzlmvl2UVmjHokYT0F2BwRJ026ZsgEceFuHEVXKzQxr7Lfsdzh8I9be9g3aUn
zXDcDZKHS71QN4Rz4LxwoBpV/rNDEZ0J1y0sFvzH4Oy6Od4TgHFRZnPWkVdlBq5O
VSig0qWCq0d83aBekuG0ATzVXUeYrO12NeTfJGiVjxzhkJPBqrlfYs6V6r9aO970
/50WrvbMCBKvmaFpmcRyIEwzmqWTEasYlSbzRjgcQ5K148wN62Txn7NqYuRpklji
XWFERquEL6A5MULDjM6jXiHSiSwEIXOyQ0bi9GM8j18shUbm7tAWJhblnGJXgKWj
YStziPpnKJMkeQKrDhmjNyF/LwCn8VivQ8nqJ5490RSqGflAHBGhegxzgjH7WTyT
8/d9CTnnkuQ1OWUESmkr+6z39QmejSH1hi/ZEd/cS2a6HpaYz+QpHca95C1QglKe
UtfyEWMu5FGYZ+09vEeid08+CbNykRkjvtZbvNmo8+3ft0WLihijpT6OzdjzxWQY
q49BcgFEMIPWXKAAFJtyc+y6WmFLDPcqZbo2ZuD30prxefZXxi8qaWboraLUoQqA
HchKRcksT/g3SgzxJ3b6ihxaTiYe6cgR4kTu/OSY73c4Bn/27W0c/UCkK9PzbNS2
eks2pSKrD7HnfjXJBhpyiKoIxjWjfmybUhfexHE8p+qf5xLAdTKfShFeLleLtrtF
0++d6HdgTS6vadtnnatSIjQ8UElWxYzfyWqi3S6VGYO5zU+eFqRraxdg7P8cORXl
7xbSbP+1sgte3zag6U2eUnHvE0GAmGdutT8SN1WNaEFkKcjZ8dtRbo71s4ckL7bA
muKvY6ZN2Nm5yhV6GojmZTxy+k8TGf6D64P4UeOqTvVtFFDh0d/QP/Rz1QxmRUNc
nG3DCLV9YnLWzALF1Q/pSmmejPUBhmVQ/W14kbBMUqeVR8tW5O444vU2xZW3KCiI
sCq7LqvixoxpsxAZtjosopegq9kXCjVu7NwyWzg3E86QtYbZ7o/rJNSkKhnsKOtY
GRWOaPIbu3HpQNOfr62EQAyFl+M3TPeEj3W15i0H7kmuHdIusSxOc0d+DBIiMkaN
aJZMq+FkT3pvJYbwSSQktrtXcp0Om+hjmWOTFu3XRErv2j8p54PeyAqJ9ARMPuBy
fxVykmfYPn/K3yr/HjD3J521T/5NZzI8D1SyHpwu9u1ZJZWY7BhFeIZC/xdi4Z3/
CeD25JgAyHeND2CI3zCp+Ht1wImpyNgJQ+J2KRcmmzfq/96z8o74HZ6FtFxSwTtu
fWBbe0idM9ogZuXGkTgPrZiWApul6CZ/E9YwXRa6Mvf5QrF56FtbGHvAwq1BwD/W
AovHIlZiazvTxWgRoyxvWPFB3ObVDd9RUR6FubocmOB+mpQR2eFhpZyXj6VI+CUH
ZA7H6NB8p61XChn64nH5DEosb/qXZbRPK1qj1FcijrJSknHaeom9NxZ6Bxo4GzXD
ixM1akJzENvAIxplW9WXFk16+HAQ6mI//tQMgx4Nt6ZHwoohqbCJxOhnsAY/x7S7
3dwkNp7mp7mFBV+DawqbU2yzT4OB+AFNMe23MD78zdfUtKdihenm9TNAOyZutohD
b45xFe/1lLIKWNdx631iqGClsA4GqKLNptVrGek+J3OWkiVN78U5JMaWS0i1msOe
jX16khuN5SvFHeBekvUeuIxbGHeJ9BYOmYKUTCW3i3uexs9mvACu+YgXHHi2Aryg
egJPqdd/p36lJIETYpNDPcu1gB5mFgTTateZCwaMoD+kkl5pT0wX5YoFpnOZXRYm
bxsZxPRfvHMDi7Q7nZNjKokmKI1vR/R6dHKtkNZRpEYiESp4SVktypGRVxp41vLN
T7m93+PAm7d7f9ntSBbFBYQ9BefqCCEVSTa59oJibumCos9C0tvThDX8gX8c5QUs
JUMuo76LhYdSEW2bavymxd0nkUZEPZ+mraUd8NPZh2tUubcBS5z7EGUfodRCyv4W
yd7yh3eGwDXxZuy9NBodCnzI7FZI2k6R32QZHXiv2VsfKloBe1SpfCuDOTbfG7Qn
1r8ZYwq5406vYtNq5mTN2kyrPwFbKkTZkq780AbGQTnkfhmmYPo6t/Q7OZ6aJlA6
TEuEAvIqmSCeaxQGSAtf3Hx8Q6+s7PALmSyn53gPbfnDD7xMB4v4XiNaxqRWPrwF
MWjsuuL5VL8ruCoCLfbB4g69eS+mszl86rQwDWORsBY67v89c9cPB74dZd/L7GCl
q/L0fwVfaZwCT/e21r6UqgIpRozp2Z6wxzPzfDDZBSPPWjmcK64F2aKOfCbDdTzE
ZnbWfvjF49w7sIZ6hnt7u2588SHg3Y6/FZ9LMTGpMs57c6y2rWsNx5stSugxeZMe
MXDbs4HyxtT5jnF8H2iVbuto3Ag3H0i4lAVq8ukpkNaWLn5ztK8Uh11NQbJ16NXP
ECXYEnrbsh3Ct9vtj7OJ/sotv7NgkLMi0wIMp3tcCdumkPKXPyU14NYpqIuAZbGl
PnITtCNM7MtsEUdrMTljbAAQrSXe4/N1jhzOiYjA/4K8qMXvuEjUxKokFzSdDary
MDF84eGa2kHUxysaxnm+rhseT50MFoj9nZgix/AHLlkdSqNUX5yAzYfT2eAsfzZh
r3zcjcj5eo28LyLDn59315q22DYDrOzEiahU7BRBFWcBjLjDTt7H78wafM1H+b7D
Y5lPU4UsxGqr6hh4SlyU+QrXRAxT9nIyu70zokRWBxiJpVbpWWbyUTW0yiyS3DAX
UA86h9lTxgdBPJpElAyfiXt6GKE8s2GOOhKkwpSmMesC48TlKdiR9rHTF2odiM5i
9P5AP0VN169egdtGHnvCB5qgoqR3fTRVEFrjjwy3vJxZYkqHTV8huxcdQ57d+Aik
6HZYb++CDM+8bwkqD/J0c+X0ZcNgfTxvCUk14uU79c2wX6QVdB5b+flKjTmf8HyV
y5rGU/MoXa5qMh59aaaK5lI2AYVK75fqoUHSmCcqqrPkPlw2ADMyu4vL5/SHj4k+
YKZWOsrD5wwF8ADCjgOXfAMX2p+4Rw2lbpUwu/bW8zqwoMMfwX5GwC25uD7k+BYN
JrTuYb5PHDGBEkBUnDMXJ9UVPuMISPm+I7Xe17uK1FN9uQnKssz+SDsWIs7vJJ+8
iEOyaRVaPF4FjRjJStvQ24epEM4HZlTwI9eV1j1wJf5ejwrPQeA/H34mGpUoBVHH
bSkgPfJhbjG41JTwokw1uwOVcejc83TPNkWmOyUVPGkXggd9G6asGna9SsLVtqHP
ZT2FuxWssQ2v34xHrLFb19wQiOc5EKXjDJJmqjy12f/3owVotkhhFSoqk73Olodt
/B37boB76tSThKcDxtQ6Tkizl8r6lrdEuHXICvK9bMtCHOxG3JkhGSfnelfOKenz
tfX4/Gn3W6OrrS5EU/f6v6bTN5Z76XCDOWbYEet1fwDH774hZGMW80t1WhqZaw9R
ZSK843kl7vKRTBeHazAu+t73PptD741SI8noIP03cvqXhcOwLRFm6aVE0oFCYJsd
zD6PjynIwVEavNGLNMdvUMulFoUy7bMC1Bjq82+xyA3PA3n+R0mmB1rYOB2Pfylc
lcKZkjB63rmaYzKMfRFPnjZhNEQPWmvwID99G9sEPRUjP1Joz0LY5dQwU23DpgIO
CheqqIywGp3D9Y06HaB/xj6sKpvxrKKyasNGJS9GV4uLa54If3P940Gycskdy7fq
R9LvNtyqvBlZqAeq526qMgpX52FoorAwciMhFlvp7GersOt0NXjGFBGK49dR3N+V
CTrHdWMkQz6v80jq11TBNj48Im3YK6eC406qXbqWYro9fm24jDYwa+3puCW2Cx5i
H7S7NSwdGKFsFGSeTHc4GrGy3JYAru3QUu6XNAkNsix0xXepMmRtXg8bZZy1S6n9
41AYuMpcCmyRYpmtYd4EklgB7mek1lJmMl6ah1+NF+QV/9ZIxgTzTl8cqnp5S8c1
fwjhmMSMeIaxJQKgLbgTfD7dbHQCzNVgIr0ifPz3Y4HgkJs5PmGmq5vlYmiKfQbL
Umx5S/dLVvunGcr5SZQIj8e2PKHQITYg62clmBSJhhSrDKnUCo9YfdZKENjB9dp0
G56eQBwhXnfLOo7CQfH9OJ47sjroayqJYv7ZCvxPdk9mqtuwdFZcoqp3V8BFY01Q
sm0u5n8v2bsRDWZnftWFLMXyR4JzF2si04lj8q7FBFRHOWfelBplKVLjkrRS5tWU
dVyXsz/BHnoKeI5pSeEqtNrwEbdAALoa9GaVVeuzPxxyScZ2HEuVSj2yWZ4oR4rA
3Trb0/wGN/JQ5qPk4ZG/GC75bwkY5Tbg/FTxqQ9pCLeTo08olmNgBHfiw1DDExMl
lDeBvGE6LWxN7yENWmS2pp3mmRdf7n6msr4LVtqPoPF4hY3gq18X+72Qe7OMY1VN
mBq+e17KJbINCbdpH8SnGPCichXjRg1Go/GsqtOc/sqEvyslU3fS2f2HQL0xm1gF
oQ9+egn6HT15nrPRaE0ojiR7nYCeJmgzoSL+obv29o0n8dq0bC1S1ko5C1cmdvHQ
TB7Xk2Lb/zfRj8dajXZftffcq1vcAwpjOipFXna6uXb0dHuAekFhnLJfNJiJNAJW
T4Vhup99BrTXZi1qyU8zqb/uEWh4TWb4JtnjOqci/oP7fDFhRdBxSmIYuPgqh27j
uKbwaFquvYCVV853ZehDQYKKsIW1p/ECgTAJLE+uOegHzrRH5DgnMMQXRVQkriYx
UEoq2Zk+HSXya/i7cuylMJ630jjmpn0xits/if71/Dtrsulie4/ZyRgJ8AmDDyDN
ZQ/xgePDg3rXcNuuNQVtClgiRHG0YMmgSblbhWIlOkF3FnqTnqGa/5z/EaCffc9u
42cGiflK9gjxg2FiyUeAv5YcJkc703lSJadV0JaXi07SX0dqOK7T0JUjqJiby5AV
rIL3djsKT2fOChGH6X6uM27i9IxeY/4SkJWr5pBJFmVLnh+UZZfDVtYwC/b2ngA/
nUPb4ay15YPhKTe1y6dmqkEqMC3q3dmc837Z6l52RKpMNLF88uQw4NGv5WSD1ILA
aakW9wicgUdASC62X03NieMiUcFVGPgdqE/2zNh1vB2zAuvIT/nyjqjixxUZvU9h
LImLOV8tuQCig6WopbHwtDGyJ9q2pcA8Gjop8fE4GMFcM7T1qPaioGWYSmfQySQZ
Pzm7L5nJYmg93k3vRF1yepveRVkvJ9aZdwC0BV7AxOibU+Ug6MWhXY+iWie1rE40
iGyoFtIL2g1b3goRAAiqEPMifLqsanqRy3xJRk86vRuCTh0eM2DRdHmUWj4nFY7i
JCnT2yEgk6xVgvBZ2KsBHspjXCUkmF6G297ZMe3oHJD1/fn5kpc6pmJlyoWhLmRE
FB3bRiHzn25QrdKvvCh+LvplXBVwZei91ClTcRWV5HFcjJL9gOzoqnjGJa0NVgpV
EfyPRN80Mcu5TGDB0a0mVo13aD+3AqQ6/F63DncWtZJqcceE87Rc0uOPvKTRKizd
fREm/sGcxU3wegmPi10rRPnpJrerY9AsaG5pPSW3dMSlPp2xPEVvg29Yprzp6HmV
xxGj2BFL6lyk1AZhx+tzYomcndOLcw3hbzapfe3V565y92jyFF7cUPhDvcmJcNUA
SobqJW8rR1cFX9KN2pppI9aMDWydvFGKj7SlLJihOyJMar3Bns3x/tHlM8d5DAS9
RR4CZxL2jY1GLvZv0m13JB9b1Nk8bzLAKYjJdD7lYpPf4YIHQVOq9+Auk2QovNGY
utNe/d458o/a9/mEQu7b/PCKn4xp/6JCyzbxoqwacipW/uWIvvbFX/xvAmyMCqQm
u9KosaOwbov/zAVg4kcH2jVIb9pamNyUVo5RpafpkQQk2Ppvrg9hiimrhvU4PBvM
b7HwXedpWVdHo3jsdlYfGKDW6Wdxgtm2nv73tFm0oqE8PlpUVEphdlt+ibzvYn9V
8pmSMI7clERYsFkCeoEj8IBa47+tHs4Ws3t/ibfGMQye0+wORtax1qD28fJ9jOQo
1FXILFrw83EQx94B9SHfdZsl0oPRbJhZ6/8M9iRHoyGEBDwuD3qLtIsOU2eShtUB
nlzAQ2JLWpC6VRi3eOdd3+n/xNFQtcuU4uCIXodid3f9YRw7wOs0t9HHq0sd2ypb
Ri673uKpKJEzhdw2Cdsw2kbCs3hQ8sbwGCsO8QWGfdzFGKz+UaHlx16A6yYe3x4f
J04To+wcmCxC/HKrsyyFD5j7/Td7pLR9uBIKobgS/13G47n9Q6Z1EZmRaCeDrQjn
GCvhFZhmovOUOvUhmj89VkypGTg0Ma2h2aI38nW2CIwwyaaDVgJ5wDKYKB9eukm1
35B7fZfvUCCg6MYHVi7STb1tdKpWFDBwJtWxy8ukYeVCnZHEvlAfNCja0uMEu3t+
y15vET5QXyakbAMfQeiwR9eZ3QJNj3TZKVcPTSPD0UrlGr8KsJgvTqwSM7LiIbwg
+N4LvEv+tDO26jJw0tus6+UTkcTZKQupvJdEdObsYtnanvOHTVNe1pF2ZZMv8YCe
J38JaMxUPavzs3/DZ/CHEvZrXInk7Ls4VZZL4hfLlFyoUbsjWrVQTzPUKxI3Rlix
OSPCEWTyqVhcgHjfa2MYs4/uVn2UvzgzxayNHA9/+TNKz5+z8rFCIKoTh5Lt1qCd
uRhCUbSMWKPbnIViHbWG0WFvrYNgc7zF/EasXX2FHdoT0ZKZ4v7P0uafAAR5cprT
tqLQTDJkdyELiZqNNgTVFSdiJPFcPh2qsu0WP7W9G/l7crMPhi/dOiTJcA/YxgzK
SYAvqmNLZttkUoq3lEKpRsmraza3AvTOX1Kf9CwPPoiApgDnWEKPKfEkVA8sE9dB
Y6duEhCmLGnZLfUn/74c7+3Wankvk4rY+6zRInzBQvbmoBbrHY9Myp2NFjBIX+Fr
HlJGamqnnVvc52CGfZtZ1keyQ2zJywqTilZ2x7O5qAXlhQ8NTERMz6mNss4nt33Y
t2ZYqJ8jFgqaLA9yA8AuK07+EVtCVNGh6TTZg3rZQK3TKHvbq4X1zFW7+UKPpNub
nc1LF/1AtknYngcn8nNKYkWK2OtVX95IhGK5znvGkntz1CNjldJq61hTKVvFg/za
7MXPxnd535jZz+oTnd6QTH22jKhMlittt+puHaewoLCr15Zm8gIZE+yFhJDG7c73
83YuLq7oo7CBFgeKZeZuXrGkWwQ9Gy5NmHcFUcCegk6bc3J0YcuYpUEWg/9vTm2T
I4tb7pk95pzsYf8SKsqLUzFaLJq7XMxtcEWRYE3lMONDw2t2kIwiQjYWSwCdIB0g
LZWuxFtQfHAM8kzoW2OS0UakO5LYtfpc4PKPC9sqdAEXTlWSSlW0c15WBvg8Jmvj
K1QZTLogVpQkZ5spamx0mbGkD4kV1hLug1rpGXKjqNS+85fyA02+vwXTXzDGoqsC
rfgTH6TJ/2VQL/tQopWClQ1KCRL6X0jU7cv5BYSu0RSONm5kJoos5lay47ALoMKm
5jcgSJ++8vdWLaglqnPI8yy/37lqRoMH4Pub1mnKXe/X1xnU8WN5QdH+2eVljGv3
w4YtuQHa+Iu8lqwGUnHQ+08r3UAYvt8qn63S3UqlaqZ1TiZv1JASenZ82Hooe3ho
CFTcTv79BQIsUxMGZ7QhHIyoZbOLZ1GjCFXv9nHHvPBfWAa2LE/Euqg8MU4pYpn6
XlbQ0FOIQPLm6TPlBFkdapWw/P1ceUBr5uCfFYVU3zryMWQywXbOzaP89f8oAkgI
spLuRjz/27BDW7zTZb0fHbDVNhxMcIqTlmai/4FBTekio1Q5pJyeGD5wK3Bvo4Fc
DsnzpIk3/mI+jnc5HpTSmodx8vnhtkB2jCwPas8xNgPXn9+E/bUih+l/fuVtqutn
9VhiaDE8rb8YDQUMVo/Vu3+nnNDH1jdZ47V55RCet9IRMCM17SyUDYVhSu4cmnDH
OT84FMa6NLa81JSNUqscM2erF37pE2nwtQqokdtBmBLgb/A2EnTTwnq9VnWsyYvN
od6LSfOnT6dbBZNaydVv5f25AM5DAvFQ6jRcRI7VGgQGKBCswF8ozo8AcpvjKMiq
6qkmbFySWniBnr7DJRUz6ywC7pEenVcRLOZ06kgujm3+pTWX+9iMtFWj0i8yqeh4
BkksRvCFAw66p5EtZFFEg91GntIGQEcVXfChRQjZOscRBIyvMjHkb6TdZFuqMOZL
a6X0iVIvHTFp8EDY2pnCduSMQyn7TsrLIfvd2Q9UejJMWzh84F7mhr2C3oquZQ8j
EXKTTCV24uBB+ZGq+NpBlo7aOdyPFTYXg6bDVVu5c3ZarM6LOFP9HEhe0W6kg8dD
f47Gb4meDyRYw+FfzbBgdi3XriQSOadgPhK/mKKPV6XMKi2IzgXodrhdXmKVrxwB
xlZV9TceMmOa8b2+RBchOLaoWzxsOI7NGcG6GuntB3+AnN9J6GQkWeMtavc54R4l
8NKgtDZbiE7VaMOcnFpXItzL56cRDeWWqOA/KHHBelj1NDqOstfsNKjlNXQQZl2V
3l+tEw/XdjacJXTVjni2wACjphQy4IUKlFT/xzggTUMIy4LjS9oObxCVMlWGMa5j
aP/qhFmHsidgSV6il8KA9Ihs6lseweYXc/Xq39nbFhnl4PCMQg7D11rqUYN6BOI+
EsXEXLTmippEqI9K7yvy9V6OREF88lsVUNsdGhWkt6TsB+kEletDBOTDAALSRoB5
TLaT3f1S4VnVL8p8DDiRQ/+w4iFQOzifYDFVb0pm1aSkAoPRY7NejmhA2X1o8rLV
yLcq4YRzvtQGavkdasapZMD+N4z2jr4tyjvoLLm+SDPP1VKu3e4FH4GmUYF+ZTyp
R+ZAH7L895p6DAkLVpbYF1YbGQdewzY9q758JgIFTiue//mGrMfUdvQ0HdtWHPXa
wgVwzZ4kODlXGBjuC1nZFXFnF0z/CfI1pEL8cSUuLh2OAAtWhWw4+HDRuE+osvkt
JPxhw7ZSM1wONRXS+mnY3Ip5LeU57tcKyHGl2bvHjk/YOa4pkwdLpqWuk5QUG8cM
/l2hPt+slrzd4XiMZsiuy1V5VfpTiZDOK8MnFP0Z15yG9RYmwe/xfcnvCspH5gZY
MsI1HNk2cAOLfmNdFmJPgPwXccGnA/hvjMrjC2NPhpbv3G+0GHO8SRCzgHrLej/2
HUjsmGxqn6fsJsUcoA2ApfPfJdVsPm9FrEKPhNK5WFewjMq+XEicYnyv64rnvifv
cy4G0Po/J3R9ORPSE6uoymNFh5m7bypD2rvHd8ki5mDGILDFrhheoMq7AK5iSjuc
+UjtabWEPB5KDqef1Qgl4FaEK14JCtYYpXyA+jEib+nYlAW76PU5ZVXT/o/ffVYp
P+w0xgh+Qyw9EkfXmE78FBKYLLfPWSuiGSshScYEcHIQfofd2SlgELjwaahYaBiZ
UpevISNmY83YjtRQB0qxLgg73hc5Sm1LrIsT0mPOv6Yhk74sMYfogS2zap7ywo1N
88T0MCH3OrefBvVy/ldkC22o3RicsU+0RlLvasJXKKjxxHLBWmLmu/LRozPCORh5
u0ZMpSbWyuLGiTg7Siy3jx8sWomZFPoa1f0XXJjaAocswKOsMPagvK4xmcEOL2S7
omQGdcUQpKTjnGLI1g+bYj1xDR6Grn7RBh6fqvXQ+HO98CpOaNxSgX3MdIzUccWi
xcI20+/P8SDtHh68DSuKoaIj9h8ifKRXmqFWj/aAj0tMLIBSQdvblcVyqA6yYy9D
t7MFxnzEGfw4E0WR7sKmX8RcqfBB01LdiV+m4IY8Vm+uQHt2EY+owLHm1y3NiN2K
6u7bFcM9ro67v1/wtP3x9yta57gSD8u1S0iPTxKWQ3xucOiJb2rhBaeHwhOP1Dij
GG6XW8ezCBhOVgtaOpjfgz07yfbHwRkBAF3PXxU3fU14MmOgCDDf6rIGkaihNS2h
tHshEDSETTQ+An5FYWNuL43MySkkQHh0IuuJ84FnNOZnVxSW8eA6VqLwMqpzX/dQ
dzIWV2mSH0OMeOpecRal83tRi0qNXEUR1whElpszxyKb/z1Wx0estdsuc9rBBQMC
HgnFtIrIGqdvw24aQuu6AmZr2DfOi34olrcMOhcIDrvbKKho7DWN2BZ3hGcSP5dK
wXh+gs2Pe+/pTC2CgNYzP4O23O5AKp0ku25NdNaSLfoA/6yMuKlvn2/fOlcelfyH
LFvRTk5gwZBPKs+Ja7UeHM4Jf6TcLc8fWAo7QyJH9wSgiomBZ9kM1Xp8V5lxn7mZ
cGFT+fErXJ0JPcQ3Bfs4hImeDtnDAoCVnGx8oiQmB/KJsoVqrwfMYV0hutKg73np
MYHeSY+STaLz8NcjK9Vr3rcNlnTnsjP4U8xgZinXllgaLIGTW6fxSPBWGOHwX1Et
0HEqWD6mNiquYqtifYm/GpxW5OJW2R3DupAT6035MzFMBqDNe8i83Vmaw+5hyBkA
4cG2WTH2E25Y2y1OuA7WtGq313VRmuCqo4pJJ2lKTa+Vl0mVYyuT/Q3Lb005HhHt
vgBwlK3sRVRjs4vjvGxfIaEbXQca1eknjjc5QBuB/4sI0K5jGNApbWXWCP5HDsPK
z+7TVIRvof05cNkQxVR90kEZulHs0YuW2v+XJW8TQvhpmZw3IBCzfHIc68kfD8qi
51AWcG7NycNcTqk/270WhD7AGz4U+Tp72R5zjakVVhfZtyu1j4yVm6vh2M+3MdXK
34WObI6djPIuRcC42+pSorOWtu2pRFSe2HUVMrWtyzTVrtYVjujRRH/nnMnJQ0Zm
vh8Ubg3EAwvsD8+vJbzEDB3zMiZ6b+RaLESBmJ49XDABt8MSvi6Lcm58PBvnBMnm
nrYOF6ssNPTtePNeQv/d43Wie0H5p7dEeE3wlRG+6qYfaf6MNWma29MVBQmwAK+T
i6sWLSRhFZU0OKxWYC2odVqpXATcmLZVAsqu8KYBS/Gtv7w3jnWZhxte833bNXaD
5lbMILDnSNSItQ0Ea35KHKAmS9B3IwuWAejpkOEcf14GSjLgxeeMX53QXwFTvYCI
ezXc/WIoBjxqcBewK9HVu9rhfzxl+rQRFTyC4hK574nJ28HblWzWV5W475zXccb/
ucQ3gH2V2d7CF1ZDwlbVIlyq1lEuUULMjxkBvVayvGQFtZHytBguWjelEk7j9dgS
mC6xd3BLt0EtCNTW7d2cbYcpBdvFZ1fDfH6J2UIxFFv4kPqkpHJ+cJV0Dt4Fnbzz
/bR6VpFHWOs2LW+eerW5ijeC2hOd/q/B/WJ4DUo4CO9KitAQLEm9aQ9WcnwX/IxR
eG05D02clEqhu0t1iC6qtn3PTgdTkA7afFiUZSN57g68cC6AM2G0jlosHXJWISnT
FcGBjjQx1WL70o2G169K2l4hCEmCuvSmP+vf54nXe05oPj8Ds+XUnqMUQhOJDd1R
gPa9TQymX5MzVN+HglNW1S7/Z3SDe4wJuP5tJ2V6/QuSVC1bg2R2mwyFWBXG/bMq
UZnv/C+Axut0Z2N8dvrhHips1kihMv2zDm3jim3ZjrrykMoBVZWx7Dhph4RQFRxu
vD5RAwiGy6PU+txs5/S9wUboYeMr0K7zbxT2Un2dVsZ3lvxHKoBqS91HpJ7jA9pT
wcGbNtZG9o2HOkptbMbfFON4Cr4cYpKgRXBgeTrtJRY3kZL8vOV47uAgxrXATHhX
aTRBofTdi/pyhXToBDe4dKn3Z7WLBncRknnnOBN1ja6xJ8NnnHhfb9aN/ED0BtFu
6xD3mVPz+Iq9ZYyzjJRmuE6bTWM4V6ljBBRIiAf2E1z9vg8S/OT55b0/ffW7yDp/
NiT4WyFrKMqkkvpIOKowi9EGKEVvzx5BBuuRJw9IcdcVckXFAPhQe37fSDWdHNt4
AfEzDwGA5nC0zjStjEPIt1Xsnz+EL4tHDMRx20yqM2gcWUDkmHwfNkDADO4pFlij
GoUldqepNdjCG99XBuG77RrSmvOmTefKTDkm+lkI4LKmLkJwtP4t7ZPBYdT2qmWg
oaR3BiqMI46j2LIQQdDUhTgpVW4l7GvHqd8wdxA4Ttu097e0knUN4HjaRDmu+NJ4
d1MKJx7E4KBT1ys11iuAmV7r8rE2HNzxIRrnH+LVjNIJ17E48h2Wdeqg4UI0wOT7
fl63g7vif78Cx9HXQK6L2OKy75+zUoSw0C7bQ93A8BmGa1VcrDDw6pQ1/6EbC862
BAtROtmJbRPJrHr4r80bg7a4sBWh+hRl66Nmf87U9owsY0CzNuLvWZI+05aByAFs
8aTxyOHqC6aaYekZrEc4Quio+mdG+dXII7fSNRbHyEPSzFhT0V874z9ruEk6WP2U
upz6WB96xMvuyVM+r9buXP8prEHL7PalUjy8bwY9hzEnpiyX/nFcjCagCXCjiqLK
MIApOANpTzxX1GhREj2QA1ZOYAi6w18+qA5yRM+07YNVjh0G3r/7Mw9lpGuR4Iq0
Y/HCyC4+atmDb8jTC9xkdu3RIUr+iWbyCdprEYYUX92BUQnXSnMFfj9XmllkKZxw
f+i/muy7QJYHcXGTu207AOG8WKg3q2kH2JsalCUnm6ouDM+Ryj4EjZMJpUIsD3fK
TbP2/7uJkpz/ip6cOY723tV2uDv08qAi3qm0K02CHUAhvPNWFf3UmPhLD0iMIUtT
+HdrW6lTksGIVS39G2szOXobmcuzgOlxykkL+OSXZev/ITQpUfEqsEu+B7Hj/Kb3
b/3tGs4akqCWjr7GOktyJtb9PF5+2PJoRfpJJTkv1ZjYhQ5mcPRubvSvdwRWmKPH
Pl0iSQxub3JONL9ydIsf4GpzYyXTrLQA9mG7fauSEUDFhjEqURzroGvg0jRoPEAO
dtIznT/K4wY/nfBLYH4mk/J5RA8iYrm428IoFpsAR+UF63iWXjpE+nezCuAVayBn
RRuP96U0DrW4+WIsVBgmEV/3U4sCFgvTxmyRX52AWd/2I1QT6fUMHlwanDSWY3iZ
SVrDOLpMaIMszZoIzWdgS/RUht1eddS/vpvQtVRrN2Z1JnR9EXRmyjYmKBjydrRD
ByVoizxtbyoNN/H8CpCn5UrZZKjU8mNJWuXsqrb2JksqBgbrCDO9gKVtlum6r9Hv
l5Xj+2N5PhOTxqx3eoQW6L3xY0TNHgAYGBxlMAlXeA0xAByWXVuT+JWMeJsN9XOa
yg/jAbTTvOrQZrDYq8ADxE2RJHIUInIgr4VfJ9Pyt+5vjuX5V4ioaOupmpYvylJq
s8fQm03fsck9Q/MICeClWKjmbeqHuMGhuZAOGGsPsNm9qUKetWvd3lkziK6MA3Cq
g5SNerg6YN+nAjV3cs+K7Oi6PTikN9IhXDVaYTWvU+cUd3qlXoRAdEFSv7mFu7i6
8seWmCxQNpVYowSDuW0NYpjRbsUV+U9ZQKmYnlVw0eiF6pkAZekAeY82STRDPIl+
LH8AUjdpgdR8lHNN2IiI5Ori9Z80j+3cyQVwv9LQxuca22htJhsjzrEdhqo5py/u
MiHOPX9iP3EnNbjIYR7KVHNx3sUTnWCfNwwyYbKyCCMgsF9r7NuAhBBjp2bAmMkp
toF/ydl/Hb5mqV2zvYl/ix45qO/JYKzWQSNyqJSc+iieCQDXqVOwfMhMDso6vfe2
pAfSOOr63j9FV06HIqaSabaS6x8+NEl/aej7WfHx68RgRVfcghzL3PcXUBroCwxV
8Or5PrpzdXdBKJVSZoCzwUTRolpmZkTeWAAiypYZ7tBzPB4+3Jq9WaZPCNWxDoSs
g/KF7fcrOa29HP6jSB6XCUv+teXX+6Lm3VtDzSzkU7Nc37ItXLloJO7k1XAK564q
E3M1IyC9JG/whiVq4XOI3XAAPtRlTyN4vppxkVjh7dl8s9EFOQaO3yEsmfVtg68A
38CJ4Qc9jLxfvb5tWUtLbCVoIyskSKnEcA73gboszFVG+Ro1ArRyy/Zw5JHnHYN8
rjTxtqxiM5FhKezjInrhjjBleMg+uij19lYwR6S/aMVDRbFCVF44IojHvAPozkKV
jWHDPyOZCakHjp+K4NvcZqz9C838Xb6xiKRkwLgr2S8ZEKaQgmLzRMkFSte9T0jl
4p4l2l9iZa/R6abyCFn3ybp4RfPsquT77WQfOeOoaoUF915g0LA3BVeTjOGcBdck
dBy7U+LAj0941GvO2fRR8OZjxryGd0JJ9im0ZawE5keJYjhIA6W/61FCtxClLmM1
P6+KdRUIBdQOZ1aAzL7pPJNdZ6JdlagdI2e7cGyDuWMPI6va0Do8p+f/JaJA+/Ba
BYWwUkd61/9hPXVvvSG4gY6kNsNAz0NGSmlaA4OMaS4xoRhUh/H42NFBxog3DpUJ
LN+4eK8Pxs+s2OHTPQItOCM7+SdsnYr0pxLk9z3qrAj5BC/tF3WiYyzyqfGkayDf
KE58aAqo7b8NRPijHEedqWU1CB5dMleA5j13ZvGph/7PfWUzC1jD9AkIm3HaKG5i
2KTo3b2Y6dzrUVKR1IqMhkzwBbXIqs8zp3C00oChandNgxkq9p0bBW4h14Q47wAY
YHm2hQ11kyC97de780GRg/N2ovWihO5VfUc17mIkduWzUabPIsFom59n9Bt1RdxD
DMQRLiA6ZWHwVOgDtCgOomo3dDQRVKR7OrXFqEGOmMynCzuNCJonqmiZbmrWl+1O
UOk239phRTem7yFJFL4hJTc0VMOvqq3S/x4uZRgTscl7YPj54PSd7bhCR6Uh6wbd
u1vsQOeF0U7ptjn6a3jLDg7WnndwkdaYpeD+qNMAY0YD9RvNyfOZRezkzbIHZdph
YLXROBKyRPrfFTvjMUgnvtZfcIIcc2Awaf0XMJ9K7TRCY50uU2t/WH6EBzF1Rpyn
WpMG88JLJHRNAQktG3CugJ3f1O9dKtzu27+/szbpkxUHkYE7Yw3SCM9H3sT3qGxt
JpN0EIxsO5oxR0SrNSiXXhH4IWDbx9PS24hRYVKFJe8oDjVcCN6Rubs40xKmwjjM
4DoO0ye/jN8HnarOL/evWXWTJVYSd/VWi8wLvrPmwOWPTWOYVYYM67FSAU2TUd9s
63aKe6hpDM6hUykyIJGAAF8W9wjVPG2sScCOq07vmGw7evh1ndafsdAMVFRiKVwy
JImYiUGyCxa0zamJlcjRRcFaKJf3tWsIn6xkyfeNuaTUvBPFUF3weMQLFRH77UyU
mOhlr3qg9VhhibRi5EDohF9m9bIqPzBzlRxu8jf1co7iOsTNHojZePJodGhuLwcg
dqFb3FYYNOICEee7zGZEKeCjOxxikjfhDn1ZlCpc16z0EeeD6zk0ZigF2Pyz2Qeg
GOe20G48wdFwd7VcNQXD9yrYANcvsoDzqgJNGCq+v2OSp4E/Jjqh0G0+3pNrSQGQ
w1+AX5jHZU0/YhiA8jic3UocCbbR/EuVGcFWL6Gyhm3TaV5wLX5Hfe1rr6q10X+j
TIp/MAmwqxob57nEhLikwhw2FMGIdg1HhkbFm/bBNi++pLlUkGTEbBh1jNTK72aX
xlTQnwbCMEh885wf5ro949OfhmGdp50yurRHuWmzuDgcXsmh/eVMBTkUlAtrhrme
ie+/4O3NexiqoUZi1AqFxM3BYROHiQnAukZ9daJC9SHRSSa52P+DrZoBRRAcnsAU
C9mUef8C7YG7FzFcsNGrxV2jdmSMnTo6xIr0Zq4enGrHqJHjU+qD07xIWq7928Ub
owgpJnLoByaiZ5/2k2cIqEysP6lTHsufsRXxDU7krO4ATE2mzWwIJBYgfRnB+v0/
3IEq9U7hQxPIJTntfExn6G5yPiOv4sZDJt5gOpZp0r/dLy6LHe20eMKup+SQCIS5
n/ZUCbCJD0F1QUd/P59hqlw9WkV3OinS1/OZrMJ8Wv8I+WNvgjJKLFF7xgPjoVxA
78jIj414qrFJkbYWZ5QYpA2xYvmCruIpfa64Z9LQ8pWHPoAmvbqnWl95mbXvfq+I
xhosBVAz9MDV0yLc4/v6COLrcvKRmbAxzdwo1+71qychlLWF1CoascHGdY/M1EUu
zJ9rmiHj9YSAUEbTZ12xWIvA1wCgTzOI16m4YEaHG3+1Pt/iK7VP4ck++xm/r322
eR8AkeNNiEBELr/x7bYtxEqNP4+QNV14nW8z3Dkak6xpEfFKE55X2fsW6evPho/P
XSxpCcf6XVAUlRs4OJU5PP3b2INRk8FwpJvpZVzIh4oTwJo999SBOLrANDiDS9uR
D/lLFO8eVtQP3byG18icyF3nhew8teIDB0Ic6yWuijTjt1Zp375kTYWci05qWPl5
Rk5OP9XRwHLl5csoVAS1Ezm33tPlq0/pZzIk5wCkBUnhBqw3lZWfTSSJEPznnx00
7N5RgA4zK3CQcLU3dFGjOcLrJ+xRKnbRIE4pzgTcJ6K735t5cZPGPvdePqjbfbd6
cmUBV6a7NAdj1940COPvPjh9xXuNSzUYELjHgTk6z+3yOU0yQsAK/uhVdZeqbUta
cltV/BkrKJLAMg8v1nJQn8+GaPqIwZ2VoEnVH2NmjRfor5hy2pyhh4TmyhbEO+hE
QExAQSyI8f/Ovoe/vivbIOfDSfTl0RaAsKhJV/s1avf28fqtnjMm1mwtvXhzbgqk
MqVWIS1xwHNt6C5XI/6iOvo1EHyPI1FmaA0fRcPvHFGaQfOVj20FIntsnVymUctG
RMaRor1v97bZP49v9NxLO7vgtHFz09uW9cBhBuR0/zliPH6xcvgSVk+ivhBI9Rko
Eg2hRhlSpO18Y6KYlCjqcSkiDtByxKft74c+f+H8TALz1mA5e7JN65fIUtEQRmmj
7wRTX+9R7wuOPUeeu6rfyXDFf3EiNHFiEsy1VngDySuPlGO/mOFSWBpCRoJEUtvn
kBLLrqHVC1EhX/eEjqzJulr1BaLvul4VypcY1ODoTFdcASi/uHOuL8yZglSjbCHF
0aTyrWHJRMbCGuWy3x85V5Y8ZCWzU6sxJ/BLeqCc3JGc8Xgsz8lQqDHZaFRX7s2r
m6vMNYY3YOUcIUXTZEGGF2aSs0PCtEtq4Nh+r9AoI+2l9TiF7tbHHQCMzywcgWdz
ZPzHEp577G56onKotEUJI90IRxzOFUs9P27lqc8QNmdxkXDy66oGx9VfNTF+0R7b
aP3ob0d6iEHirM/JcMBvKRuhZMRxceHYkb9hHDK7hKj0JG6ibIIKs2ycw/NU7KLe
pwokLQusJ0OgJt3Z9VGFOeRt2TaZKIWQtex+Bxj9z61TkJI0iVxIaHiEClxk8lN2
hckCWO/ePun2TDBtdJT92mefTPgCNkNU6RuCwVEhUYGMOQla4LpWpPhUeTC7d7Mb
ucIxvGXxVDSqDXMJgqHtNUSfLijHtyZCk6i/mrJ1Lo+Hf3MLq6rmHIJ9lsrBQiJx
ITeknQWHjnwYChrb3jtEQ8iysPqSmRPLhSKKbbLZ2uznh/uv/Uf9zrmaJbTZB+Eq
+AUJWB2fsrUbqm5Psv3AEF3unW1grAlnMCVD2TJVA1k=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
naQ2YVN70Km8TaWx3g8a0Ngtl7nLsrvjwjKRqccADNvQpBF7m6kmzWF6cMyQo4V/
676JL7bMuUrh0aRCJ1qLveBOQbTHk4XVa2cqU4FOasVFABujxHeif5qYkD+3C5O/
qCTJlZhUNE1MMHzLiOMxKO4N3aebpYxJyC0ylkUW8h2vRWYdMh24fHFZuG6EOSEl
dnSDjwW08lddLmvbnxzS0VowEXs7SjbUWuJZnnwOQ372+BC3e76/nlb+jAwWZBfk
ALY/Aj/29buT4EV3GnG44KBHk1k3zGmPlyyoBZgD1OqUASxqSRHHYAkB6G/+UT0M
0dYwIPlQ03B1bObJgMDwdA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 544 )
`pragma protect data_block
QBX+DRmMMsYdBiOklb8WGp4OJpcIe662G7SS8I0uMqDHlZOHJnfM8v2ZnFm9sTu9
x7xarzY4LQs/hyrB6LmU0hB5EAXpponLRoYZ5cIlO3nSc1P+cWIbSoTq/H1/nk9p
Rgj3wCqjVg//CiFl8uzlumi9E3HokHdp36u72YXvjsccVik0CuBf6JHsCYXD3ELN
48KMkE53HT1hAwO64JGiTOa8wezhbVXyP3mXbB8+/gpPc9Zx0TWK6qlXtyl5E+jB
ZPul+9yxlMeC+ni0PzfO8zTBQqeC/s7DVD7NH/dhf3vgftiUaf4VtAuNsyxM5UWB
+4c3sn2DiEi4mZ7Ksg9tYkwEMOIsXS4uchbFKopO7s5gAjL+QAo9HgGmEs6rf2YG
JDyKlpi9sFKveXJTCDkqvd6VwZu8oTJq2ATU+ZkrQwkPaZAxq7fNCq0e5S9ETj7N
EgPOGfqEdX+8SJQbDc9qpVjOyqoZJv/AZ7Mcz7OjWglNoACJxRtNImrhntnzvB7Z
k9fZd8mGBy9pQJ7brH2Hk//7c/pk4zYv3MPO2MReMPJkUu/hz3V8Y/a4APV1Zooh
PZ0Oh1j1BoGMNyPCt09fFBLmDvJxCT1H42iVEfbNOih3WIxlYQ9QxSOMDEBwkL+Q
eF3mD2Kae2kjv5VFh8Bbo5JWgqebBqiSqClFN+j3K4jslXjMxVvjT6difKUlGzzc
6QVJTd63cuxrJgtfYItb3Q==
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XmBKGxIXaZH6kKRRTAkQ4M+mnqYL8lTa5SHKmymRJPlJwDP26hsRpTPvYVhSx2DW
+Bz+8ixdZ/kY8QL7W9ttuEyz1RhuPRDU8OaWVH8Kw5fQjYGk8tParVOsyZVnK+k4
erfjwYpPPqtuK/nspC3YUiUke7lwErz1EM/Km+78mNQ6fblVhogmgHIHzGsMtJdn
ohP6tJrmV85m6TbOkpeAkG859RX3uLAArtVh4/Vz2w7dD0vmnF5AUsYfHoJIEDIS
wFGtcljEpBpyBuaJKudMafayoG8iSAC635O58irKxRija8ps/kDMkXnSjQrDvkaj
p4zza6hu/CsxP9lSmAtXtQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
ewVu/hy1aPmEIsohUpbcbLZuJPvljCSJk3S0OiruAqZE7AuqOQnJgXD1p8qI04d+
3IMzj4Tj+39A+Vo12miIfBzvF/0k58yHZy7dmA6J22PBUF7tTJT+WbKNhDppO5vq
LtyBkEjQf5KS+ZKvoYHOI1dCJgmJ00AIUdwhEAeuCPtagErN6yrU1+2aR6ay2fIG
i0GsQ1+qhdzEN5MTCmFDhCZePFkj1aF+ZyMHEdiQ76+/t3SQFyigpgWpazn/SQCB
csFcrTveWquordymL72LDPrnn76U+41npkebeQ4O6Ffa+HALwb1rHuFKSvzBBUYR
/xC/iOVWDtlqQBBiuojSGvFlZ5nyIb1nV8c348w7F50biqjjH9fAolYT1QkZigMt
De9UAuRb8RQn0kY5ZVMBJWu2I7FT1Ho5EeDli6L3MYoDAoRmW+ieUCvHysWpcd2R
RqFEcMNIl3KdoyF64jrbmq4zVRk8q0725iO5gS4vNA5AfvYk2TnN9S5qBeUoIXLx
Bie4/p8ayG9af2FP/K3ps6u3emZyNu0a/zMzXblvhdVhUWkKiwkEU0SSyLlWUEJL
vBio4M741tjvbrR05MhOeEDirKJ6HHYauXVKvRfnOq8WUN0cAkvPVI3FS41kLfhn
93kqWyf5FskyxPwRHjVyBXpIjXj0Iwf+lkhNgRzFqqSep/EuBYtqRtb6MYHAxPGj
VaZuh6e6xrYRcIzf3SKMw1iCLREgKm3vy1gqCRU/hvsfug1gYT1+NY6n3Agf2WoH
Zew3ghAH4Rs9XMfPFKJbVKMEzRrCsCk/jsmRrkJpPx8NT5keNlulbeWBN/gszHSb
BsWouTKwU2utHBgn2hzK03BCgnqFFw6z8LVV1nubZT61AQkJySRhsf80djgvCVpI
6FuJMtwCMH3IQyZ7KDmWZcvh3PW2xkHWbD5OIRZlnhc=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RK5bMEgvLMmpxORbFf8VeVV0e0gTSKQ0mf0BSJQ5HmCDtnwWOtkkEY9Z5eUC0U9m
T8WnvE0cheLFDPsH+2slnImujZA5bJ89PTFDhOBVRXtuZkKIRGqMfulBDGWVzc8G
JxZdDKLrhyztUo2FVabyptO5kjBUggtrMJQBI8uhNmcxWdzGsUkWqOICyWLJetVY
Am+bpCfIbj0+AkOYOyXZKq70XTbSWqjf3+gNT2RyEIZzlMUtx1ba/iNa3wJ10Fpz
UcbI2c5i6HKtjl9tGA/aQCcTE+41snJWsKfXG+hN0F1z+EmYZhn8tkZ3HP2cyWcO
ZSBmkxBQe4baq3g1AO4qAw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
yyGSEDzSX3kfEMkhflw7uhvZOhE7QYA1JxQPgCv9ejvxopCoxmYFxKj7Hb/CpOrn
C7Xk4dkghzDSzGO2ZgBrT4J10QhLQYL4eUJCu4hNE5I9VGDrNEBySMYn4Qz6Xaf8
pLySKFRzNllymD/Iq5AH8Bl2UKZcBT3bSwpFHmEpeb3vVV2PWrfkm7YqtG6gNHgd
kmUYRnRcJpfmjC6LUmJsIPEYk/DE7K642IZ7YIAKxQ5bwr+coRHJ+YMAFxiDjk/L
4l6kfyv5NyKFkiSsv9raedMOWVQ39ozADeKmWIjpriWKn8qqaV4bh95rDoOBMbBA
8Sxx/XWF30kXXw8t9EAD2ujF++IYgpNEyok9sCEJW486sdb3AbzID3/mhWt/Y8CT
sIkmDcOKYCmHEOhzSLcQHyWhirBWpnu/7cYIMImFggW+9zxTIWKXi9DjtA9ETQPZ
HqFR+dWQiUXvsnn4UYieM0SGzQBkRZTb+ad4DuO6VQga1EUDYRFr9WMKCEWVQ65j
zO0+Qmb3ZZObTEDu6lvhJixnystm0dljSGTwAvhKmFS3lrD3X+5aZnsMF5CRGMwZ
P8B7QVEhLmbwIVUYNkcIym9RNp72rMV4iJ4YHUmeBxOnrC2oWkc5X8IHKun7ctjO
3S8G6ujrAkHBS4/nsYGZH5rn/ZCrMNSxqnHJUG6pM833dOzI/5RfXnZYmEfWX9zw
pW0Evonw1jIY652+eA5H901wygts0ytMRWglLZoZpZBiS8ZmUkJ1doTJynvr+eFy
xR9nFlnQcuqE6LGJ9rvwHtQPGUda9JIxZcDLv3+jeNgOovGvz/9CIL+k6dSMOFy8
rw4nlDiLs3l5eGEIMQmT8YyxpmqFoA1+9w7Xqvfvi7n6aEAsFyxDQl5t+zSfMTvo
blJuDzlBd3+fRqMt+wi5gUMtxw+g1XAAtOz2t1t+Fj2kEiR3+skgByiLwx8y5ykP
Inv9OshHLzJai5oEj4S16Ztno+nKBQn6vxuZ2hvEuHUFWe5Zl+dOiLHUneCLzI2E
DypjM1B+oaWMZXFS/h/0KXhhZLjjATN9C59RbTQ7tJ1olsGVB8ZGkL+t/G/DgZYH
TZQ65pu87zyf/V+v+/vWWOMXMX3Hz8bLrJ0Zd6v7bPcIJlfE5c4Gy9zHYQ30PXBl
J7OGLFdQT9E0wpgUZfGaA2rGtmlSqkv23l4snaXLpxkrN1WTlfCrgenhG+KbhVn3
f4n/f+x+44O724IpEgARLSbtqEFXvh3tF58stKFRxcl7UoL5yIZcLnr70jedkK+z
RjprL3bcRyVjfupCycubesqllMtx4rcL5ZJiKRhUD83ea5PUqfi2aJe736oAr8MB
V/rN1hLJNRoXIMcyR+C7PMmDjduBYazEQsNNo4Iy485ixVSJ8xlMRQSZaOoSGx7G
Q2oO+x5BF28MbC0Keyg9lWD1nMrtIK+CFhTHtotKKcs21Bw5QZZSnD7Acf1TfSNL
cqK6T8knEaAefI+aZRXHJs6ifOxGBRyA2OJj1tvN93nccSaiQiIhGelqYCWoAiEj
lUpMHOkHcSdOuH9n7CDoV2SfQxz/3R51AFSJDpfb36/zKMyI/1o9G2d3j8ODpseB
86ne8NOCRoVTtOoQsWH6vpg2SmCcwtM/jZzX/0/Ln/PFV9BOBVq9rMNfvtHKAF/v
eP0kO5guQVW2orcu/YVRzdA+C117FRapTKSAzhC/s5HcckgT31AZprypZzaax5jo
e6+YeVI4GBvyyvWd5zh95lo90XoOf2Lmb3hL3hAEZ1RsgjvtK8gTzMHwAlE70Ecc
0vjwCusWXl5QUf2icr9uL92n25M2/vfiAa6rPNC+IWFi5aods6ouWX+QHL7aiYHl
5HGeMK1tN4U7sauu4F2bPOiLvO+c0yROcmkGM6bqAP3dKGVPLvJ40OsjMDkKs2ba
h9K8utxqxZV3ONgHHQUIShO4voaoO0jGOL/n/XEV0RziryxgDCiS7aN5a1By8ZkE
DC6aqV0fGNC6DIbQn81p4dC4W+pSYLP8uYH6E5d1smr3vh3wA2S8mjrG98tCvOwy
XvIkLuYieiEu+X/HvURaKKqdB1LkZ4bTPYTMbcir7t39ZK+VuQY0T0ZbTr8CCptO
6CNz9uY67B8rzrYlaAtpKhOB0SmKSQCnbbFnrGq2YYnl+k7QEZbw6qBIBUTGuOqb
QW37ahOFc1MumpMeTl/XLuRV2IjBDP8E6eUy/0dmc12quqAN6xzLq+ytBMBQ2kEM
OhAByhwbOKNX6E/54lz7ZZW39u6C9Q0iVuU7QRrd1D4iScYTOaE8piBG3ieE8CLQ
A515xuaYCRo8WmGXoSTLlDp9imtg28ZKsxQNQpdvEUgasB394TcM94GZJg8ZbnZb
hzD4owabEiOsgaS6RYkEHvThKIMYMnOf0NfioxKejRQYXdjmfV5modshFnsLymzw
iewlXBygJsV0HnqUm4e9irVlnOKZr3w3zfvbUcB8JbRFm8wd76Gk6cQtQB0csOHG
E0YE3eEkIITlCp8SBtbmfJCf6LoP9997WXk7Rj4UeZK9/G0/d6MoE6ha2g1rNvGz
nHDx0mxikgmrHyaBfinsm1yklDsMk8U2mbu1HIkl8c0cc1s1MCPP+Zi9aBdCwAiq
pQPGfin+TkMhiGZ7I9LWF29R56g6MlOHSxdOtN4t71k+0V7trQi424J9YMihS6Da
ztAftIUYCu4tOkjZG/RZQmCGmnwJukynAtOMAGDBbmpH7SyoEKQggaruU4+/UuWq
eJd67SL/0T9+JrzSq1BX5zaFF8Tvrj3iImzybOlCNUH74kXJECkpKaufm+Cg2y4k
NQ9JxrSC1tkYL5KgEvcPnL58ZRFDos3jKzarjQwZPZflSB531WitoP4m+aDK5vGl
h2uuTP41AKILNY3DnuIqA5/S4Xv84g3NapRr2gXHpsOUc5YNo9fI1qNVsrYYZTLo
MimFpH6eUpaHmWRJ6YcPgKganDO4cSP7x6b3n1QI+9ph2RGRZiNN56gRpQ/aRt5a
lnG96gjwbWNyVoq7V3ZlnuwcQvbfgbBrH1q0X5HH+afg1TO+GH0RJqEWNoXRuHYk
8gVvHt4bBqtF2BxmnODpKMIt2qfdjjhYMHmdflALvPxz4PBPgOgMxTy2ZKQSPmtg
YfP9zbxoOTOPPAWl4nQ7wGpdE1yM0ukcHw5C/4gzlNjZkrJUkc7bPPZP4LDfH6PB
/vVrSw6mHs17ShoI0/XDKHao9HvaxET2s8siO8yjiwTMK6kwlzH6itnp2hBjGe6s
TyyxGcoOWZGJq0zf0PZRWdomcUewrPnj7xgUwv/2f7EK77W/nDVhsi5nS/4opOfU
rjFIuLKUaribyF5aMNq4gjJaBWxzqgVUyp3Vp4PTi0wETi6bCF/G/I4GPaDvkb1V
i99Fqj4H7/WHrfTzwzhsZ6pHAz4vDqPCYOvNg7GjJzytpZCfkOPitJ2Bt4tnD6S7
1WkNUkewzwqPO3qIy4g4gygo6e/e+6OIadTVVeD8Q3o9qAP/0bAUNSQHvKhj+7ZG
Y3r8DDA7qAScrzwh6yI9xDgjjpyl8PABl/lMRb8gCopkzVcFEwWo4pqzIl41yeBE
Bl7v2/n7AlIZHuL718gfZLff5EAyiyvYJ72NT28hgj8+dfhaZQN5IsuVx1WW5uTk
QPYz8vcRs/7HLWY3/rthR28TW5Z39lI7qlu3rXW8/ZmF7ZeWUTGHAnZJRJ6wxVPo
UnEyhHdN/GxIa/j7d2XiFzDvVt43/62VAj+OoIlgXR9mjjAjDmo1E1e84HPjvLt5
fA9IXf3j4o4am1zrqXK+7rwPe3wMFhmIuzavzGqVeyBrdlLi2L/oXk8fzBw+8Ooz
EqL2ipF6GVzfuLNhyDgz+w7gnKAlC/Z8xvirS2p9PCWOF8gdIMxf+G9tycSKtrgn
Q6O94lzNBOjqXl2zEJtxpPYa0MvAKEN1CQvgJWVjwnjb1IiznPbmtj/sfSyxXRu0
prUtXajAx2Srlrh7BOVTZpYdgLfhQa9KhImaWYuL5PEXWChs62NoNkZmsf5UC0Xo
XZajui5BFtA+fGg064xXJuvDwFFzERiSKSNExcimDAWCmwZiQ2n8zuqwvtCfCFUm
W0R7za3T7pHrpQdChF2QvnAY9GidihBBXEIJAAykLa379kNkv5lrH32NP9v/YFuT
PotCVyah9xAbWnYBuVM7YABK68xWkujGqgPUOJh4NHdNa899hP3iwiYUUPuCNXuQ
3YTgwfxXOHZcqTwacm251IxOyGwIUEAkqLllZvYWm6FBCGrWA4WCWWWH81V1ktck
dL3JnH2K0R949v/7JXlXNRj+kaZkNiIq7LIIUBFt3xBSnhsvbnOVMJLa4cPjGpnm
mXajoDUIKZoF2FxmWq75Z6k0Mqi3i9/lavR+wImRy4JGfgwsSs9N50XGBJ6PfcEm
Mutd2x5wXzjctyJTSsKjzPpQ2+mU82OiSJIgPtU8lMrPNyRuJDKwPHl75fXXS/ZL
osh5WCyGPPwIF4qiUgfMHnjsgwblKImNMDSM0rRJozOM1Y/SfJTSMe35Rvs64w5P
C5aFWVMp/OTUmy66N+Y/SAc/Fhi+ogy7+/g9Rysj8oPB2EltogjjORmajJttzl3P
9jLKaMaznastEmvVhg9clOtXQ9bZvxk47Wa4e/moFx3Dil/4XfLVP0QB6xDszPU6
nqxF4W24gqZVwzYoOMfoY7+wAw5Ds07iNJoRBZ4ip0BH5PpKaewiNNaZ42t6n8p8
3QZ9TjllPR9yfwZKST6DZFomtYnhQv00gIL4R7zC7pai9BXk8mA8OnFKO/UFn3Ke
9F8Vydr+xU5AA+w7QCoLExIObcoNL/bhYJ+UEn+zkYILnwDF8/0+s0nK7V4sYYnk
Nxp+EEIajv2LscSNL2UrJ8GzXdPHE11edqAFQarc2fENNUHqzZlP3xSkpT5nKJrI
8VACvxm9rVKIVKvKCfM8i3oAhjauVjXkWzLM7YzqiPDWGMFCV91sfJC0DTYz7qMY
ROX84Jz+rbbnY8Q1QedhUFXYYC44jhdw1fwO0BGhriMCrLPgJQX/T0Bit30E6FYO
ZRj3jN4P5nTWxlEmAGEbgWS2QhWsC+1oM3wFk/AC3d9EvZ/t9K/IGRPnuXTeh7fG
CA1Bi8yepEXDGsnSw7BqAopSdIYZpG9e4p++0l5BgobKHourHjIey+KXx1nXOdUz
3xZLhhPl3P1k8BY/OfYDbaz6fGx/gr0V8osxbXsSZBlsCsbvma/3v+tVnmov2e4t
t5lLTt9u9nAj05AzsOSndbwXZNhG4pyOqCgon5J4i/coqtKFDNoEjwEzCY1ncg4q
X4noX73t5nJo92mdgdINuzLZYaKTOjCBQJOFgXk3h/3GjOD9yMOF4Mxn++zyI1eW
JZdoKh7QvYyM3QqOD7UNZaFqxQWL9KqV7uaggNC2b2QmOyPbYeWt0QJGcLO13xL8
aACmeg9oyYW4zQiTGx501bfbH0YcJMu3n+hP/DcvV/fMnnT3sJsToUp4VojTpdMK
2xVWc+6oRzFAz1s7hSxyPdzx6zajny9sWmaeIVos8ziNIt4VBLu1d5q/jBXinPzv
CjWP2lmFcH4bwpY2p7C6tjd71MUd6wvje1zHcgU+T2NI+koL9sw3WWYCFbzwo8wo
s5TG2eK3t7AWzfXwRrwHOUd5MnbQuuW3zU1j1rXg3eM8VHG6Nv8WWOWLqCBvbUf5
UKPSxbS59jMSm9cWR05pf2nNXtCkgk0uhncMo5Pa56rhQknuQes4hp7VJXEKOSsm
MyMsEBIvtNDG7q6QxOOXH5Eb1hqtNQqn3jj9gDbQWpChxdzYMPTEF2iSFLBHbgqT
WaPty4A4WyuW66ggsmihHhNSmEXNEzOfqpMvT0iEJgwBMtJ33HK/HYiVDUQXkJqo
duaEtB6KhxxKj1VVVO28xH1O5IyWaVcDhkA+HU5/WSLyS8FIvsZZ3oVSp2kpm7qO
KnMcmxSo9G6+PUtrkGUMUmh7lQE7eTE4OY6tcAr2Zm4wYe180vo6h0Tt+0go5bJ1
5FMMzuXPPSf6g8PYe/Y1qnheZd//aBcQ7HzoC79Ms5ZOEi9G6fDykyGhpzuiVCGI
2g77ghIz04KaLbtpcxLR5q+xWIvn/QO/jsw3guU+GED08sUK8ltFBbIGhOTX1X4Q
AEz0y6hv3y+JfDi4ksJB0upZGlktSfkJ5CNSh/hUjoKQ5wPmuMruCEDe8MWWDC3y
uyU5AIcmkN64iUMVi2gJV5u9edhk62li2AqJmShwNXPvgMInYbawbuB8yNMGqeZQ
EJtOU/Uc7fyCbk23pNZtdbw1N6zjOWPvm3ExjHxoM31l9YW0dg/KI4JsYBTl9rMv
RWGIP5PN0fcyq/TljsCR7UI2uYcyPQJD+lviyVIPr9butiuoonEepOWuGVXd8TSM
0I8uvQl21ctFRSREqmgMqLVRZM0UdQtMjVJT2X3RWLiKUOt+A1zIv1htJ1yl7Ooq
HJpqukvYDCYyVcxCQ/eYWnXguEPTVkJmhuocmRThvVgHh110/sjx1Jl2TQpldlMz
cNJcOa3d4kKXUJUfemXiHQB0weJAYhCXJjiQWjcO71cf+WrK3IJvDQ1bUHUXL58Z
xMk2442wchbkJ+nbKQwFCaUkNwUy9dvcNSmT/EOeyUT2YjP0T2KoOByW7LLArYX8
e/OAlQBu5Yp83QUNDFHWdinYr5uK2E13fi4ueyyCGTTLn3Vl82AK6j3nl1iBp/c0
IMM450MEsCSr8ZZeUlY9GnBeYL6gBqUdCKD9LlG2PXxE7uDSdsJoDaW2rvvP97JA
2miDeSUMZik7VIKHEpWuBMB2LvsS2DRj3uNeb4mkE2giB9lNmPlegS+yNDzg3JLS
xCRYwDOXQlTYtURGI6pj6Wze3GjeWjDW0SuZsIweAZz1MDWyT/ww6QQLHfBOS6an
Hh7MLOATzklxTG73d6VSbcMCIuHGX4nyPga/jWK+REbgiKxZVaRFbVINUPORT1mc
i+pEYCGVBLElovwJftLwutugTt3qIr9vUkNLy3Rg0jF0VrH1EYS+drNMTc4cP2XT
fBX1jG4W2JszxYUelx9VEXdwLy6UnvRFg9k8houeyn4y4fQCcsgkQTg1SnEUy945
Z9Og/bKbQJFk4/+2+85plgoSbzMfaPOlGRnqmVFqmD2wx7aEWXucXZRrYXbuJPZ+
V3kmiOUm+ujxA8kvTNfJgoZLofJdXyyz1efM1VQbPRf5HXdPin/TRQ4jlR9i0fG+
01Ir1zCXyrgvVXPk2TwRbqBMciQAgNCjHveXqK82Z9rnUzlF9tcOs3Qko0L/3Ul2
PB+zknOpUSlKFzA3HELOzMllwSECXPFjIG3liA31g0qUc6n5LHTEOa7ieMc/phf2
oUWpHsSQtHSESSZAQL0ouuYMn8sxqWp4Rnwo1VY0lHiA3ZAQ4Z6j6XqDMFDLfEWt
u173Aq+NUNGj7ZO8HKzjP/xMp3YxrzItZW7p3+Q2MwF7U8/Not19J6BkuTgW9+6e
gRagYRtG+Pb56ebqAmc7LhZjyWjLlz5JH4NCNZwlzH4YtPePXFEN8350CLu2tg1q
3Gn0CIhEms8ikuecyvxLyO5r5i6YJYc076jn5kkqotEpwkQshxcMExh7W/v6Db7J
EcCAgq+w/wOw6xGJVW59HplUrco5vki5P8Iw22yqfJO8KH54Y60CCmVuhLgOp2wT
6sZKLz8gS9tp8ELhEhgjJleoh35cpP5Ise2QiTE4GCbcWZTCe0bxaLn1l6GyMIMW
JNp4nzSBo/+3KZQeYfKWHM4Eb85jC4u0XtBILhC1D9Wg5HR6BNJ78VI8GzMBlXJn
SPo7qpF5rT69zpCsbSV84jFlIQIMuAo8w6ICHiTbB+LGVIE7mH0EHZo6HZzpHkUl
0mXRdrUbnE4IXV05/KMc6gehXF2xFwJKPUxDG7TgwXToddfebyWfjBYlkCIIhwz2
6Ge9KSu8jD5aGS1AvSrqHOaUpGzUQyyeqEyttipgocehCe0i4r0IHDpn356I8Y+p
PdSsvsV+VbqOw87VazirUzzx/aQYnJou9AAhXhzLFACtVRKxl4NrplBGY13rbXm2
VrbNQTGrvfI6OnYByavx2V+s7B3IK9/hqNGmuzImtEQNB2qI/jdD5oEGAiPfI0Gr
Pttd6zKbbH22K3kgC1UuCqZyvPGq7I0k5Zc2sHXGZ0k/lEsz2bDobN84k93w2yii
F2zPz0s+DvKhVavDQ/iphCRUn35HeRos9HUOaUfyWW5j2lDnxFnks2otA5mOACns
MeGKa7yX7IAsy2MrehEfhYLEh56sPoWTgQKhVR4fHMBjv67lhK3uNJ7Od2HwcXvW
Goo8QwDgGjl8kBhZKRXcNwN3dWpkbQ+RRYDjU+5KUbfPQOpF8rgsK20ssXPI5ORJ
ufpME31uFZIUVRSnkc62QPPK4r+qb7ZaSJlXvgMfFxeF/f1w74X7n1NFpOyB6dSU
DigKvB9pDzLndGh5W5SKsXgHFhFth+lE+sIQkXG07YHh5ehtPRnRzKf5aTkxP7se
2ofcLkwELNzf/e0SImsIMRCNh2c2vGYugDLdUFErXqsW01fGgMuo6q3RpF9AmzEu
CA/a7175fylAtFzhkvMorBDNrSkUK8JtKnE3W4OmSb45Z7IEOiZOAAJEQKF9isvS
knRufo3qS5Kwqoy9gLWy45Jr93Uy3Ax7ssPlDooT15WyxV5TJQMnLWz1yBLlJFbu
one2SuVpQdnCjT3ep8yLtAyCFoM3xhrUdJmxECj+qSiSN7D/1DPwp1E+i+kMefpG
YwW7WwgANrIYoR7xixbyPPe8LXd5Nfb1b2Uv0lY3dTT8Uxo2tf2Cwckfc1OCKe3e
NtK6N4kxus92HrohMoBUhxWx1jd+QSW7rcb1eNT+vI3eNL3Pvd11GBbzmEl1nzSI
OoTaZphrTp2BScUhaeEwDeIdT4rpQEU61hP+VD0J9NM/n9FealtpFJXjWGVb6Gh9
TSOnJFCLioVprj2QN/8a4IbKZvULqweuaJHcZ5/zMef1hE2NCyKEwGY1xoKL7TRk
vK3R9FbtvDnQjpbEyUy7Ub56lhq3Ypi6coPZsNRSI88WGaTbmKRAsHBH2QpcKKkC
KQTujXrfmBOx3kJ1YJnC7SlF+Be9CRQVDxku0d0F8kUMvkM4qPc+uXYv4xxIMI/8
1CSInaSIhCyfT1zay0XHy/x9jph2DW3MFfkFIDhPzzhuJRF2NJ0Q+b6JK33wt0W8
8N4tTsriZTzE82iD0CVJCh7gnmN2+60A/rIkahhUmx+YolFLmstdwQX3x+0UNLTD
pAtCYSQLjfHAcR/kUqC0bMdVP326QYp1alkGjilU00a0l4Pdb1NkayC1+i11x9Ub
imgdfGt7FqV6tkBXl5wlgIZeAY67Y94/e2GnQTzosHeg0IkM0XLsEfP3Fq3tn5/k
z35yGAVpj7dSu73zd4XtXIETLatcPS7+kE8IYIDeKICFnEeaGbiVpiZL5V+b38I3
CExIIxfMKp3DGK1m8oSkesJV7ZthqOuiD07WTgJmrZt63O0WEnVPXgUijsxKmbN0
P29Ao+T5n7F31GbTn4xHHYVuZRpHdE1OAZNXOrMwdbd9fMt1Bp8ksa0ix1gwPbfw
TE7IIqJ7BU1aKJGhyKbLF6QPeBvfBbx9y00xiyvHAQNRMQhTBcMlPyatahOh9Ma5
Na+O9MBF7WJKySsmLzDGyR0QBpxiSgo5Ba7IZ4nW/x06nBaRkx8D3dD9aB0dfo/i
DyyX0GJAzB3a6nEomhuzzWTSxJhl71gtaw5avZ+eQeRCgs6lFTGqmnfyrU/1idTV
5+RgHVM6ehfILqWzgoeyiI/52u6N0d2MCWtahRwkaxh2Cg8EOIXcq+GHrJJJIZGn
PRFSQ1NyygWw9S4j5LgyNMegS9OjqPcymbWXL+Q2i4Gg600keCqWq47RddJX3d1d
lPtshqb/Zb+xOG7SBnXWOIcJv4veRWzHs6BdnHlHkB/39jgbst1cpA6dlxtTTjDC
6PWbtM18UgQrnDJk8FZzeMnjNSC/ZAhB4QMV9IGYF3EAlhGpwHHNhdWl4xWZCz0e
lHyHvi7YfbQxtVnJ37T3fcEdzTyf1UuC6XgDbPw9riCkg2Q9H/h/UG5Po0xFgn7c
iWzWd24x2FaLn7a9BZdwwwY2BcdzDBWbxGy4LKihhbtaopidyFBnrwwjXg3KV8km
qNhnbk8gfuZqWTAA2pfOzIo3/NOdDbVPv3bti72aphYvEl3Zl1wdu6VVNT81XRcc
dAFogu00NZK5sr7BWSfMLCHqBYIS2DfNay3mJoruTYyAPvB3b0V+zjg3huPu5pPP
eqZKXfDvivyOzCeHh5ONJSCXXwUJQUOCYZEPoHKPDy6JxVj0oZEAUR3lqShrPOhi
zWQOAXZAU2pasNMqJ7D5aLyXc//Pb3yN4ipPww5FP8SBsCCnkGgGABlMvh3rIV1l
qvbGp3jA4JBGfCxr6V6Htmxh82lBed7vhSjS20FELyahdR/cQ1do7jwGlxa6ep/T
oktlL8qYvllcIQa8rht5O8dnmrNSCiqdm/ZBpBPm25E9uZoFMZYWSidMu2bd9oEf
NmrGsr1YVvZfE5xqI8iCRf3AKQeqvwy/V9QBsNiBd9yJh5WRBCIc3uOpPRtGKScL
/YQ8LpUA/EIF6UZv+YTIh0N7plLwQjCKCRZcuGf7eNS9W4e7dUPZIVhIpEzpL7bL
thjc389oEZrvR+slKOZt3kWlSvY72rBg1HyEHbHfWCY5kWHx0fRsa8nG6K+sHn+K
8fBZ0iBQ/4NX736au/aGjrUadQgp8jt458Q6Km7lozyG1ZrjrGbMArVQOvG0TJET
7stxa6XST225YJSe+nY1z9NNa4k3k6mmjesX1UkbSelER2FCLiTkUffKXpJnkHDn
qhRglh+9/zUb2/pbhSlEJQK6LP2IR654ELzDW5BQE++Ri7k+1/Lul0yikKvWwsyg
JRUnSzvoPdgkGZKRNIHAeEaoZxQBPpj4P9jnHEcO0Z2zaRCLFWqymzDjQswDI76g
hIhUjZJHyr0rSbzlFllYAHx4eXDPCCX+l5NSA4H2ZMR+w60b9EwkgEEjC/ByFuNk
3rDpVi64G1Ltpal3c3swwiznV7gAG/qo3f1trlByNQ5kIQKRPfaJTcLa50/sP9GK
ajXj16DBbzyn2s0DfVnaEm+flNn9+P/585xArMWLN/6JfUpfEUdyjMceiC/g8iwv
bIXouzsfvfhrHGQdko+bKS5RZHBn9J2BoPy9PAnV8bdSCJ2h3+QHZPyVQlAESX7D
tIQIMo4uTu/civPv8qk3eQvc2vXHqx4eaVTbrMMifGjwk3gY+Rzp1XMVOouwGmQK
W7CkQY2VdURry8sAX77p47AhJk5Q7fuefwIHOuSQlG+bnVtN4VZZcQpBnS9hqCqZ
JNK6Aegbt4VpH1mxSnGNjA4EF4yl3xl8ryrqX8OP63P50q5FHeezXghrp4S/YU9G
YQyWRPJxnS4PPvkf9eDSrUBbo+ud9zEkvi5l6r2rcy/NuRde9vLwU1fr3hMqz4a0
ppMwBkFcgeHQRLM72mHgExhHJTeOstsCYm6mQEwqStW6lOu8Hka0xTf9ckCFQ7hT
mQ6f1qzweV/M7hTAg4ipAIKBRBcRNTyFhAgnWuEcPPIcixbWlGFfLS0Uhdqj5mQ/
m29SM7Hy09P9MGsWltTYU0I3vIrWAjEzSEmrGWpYa0U9gf1P+s8ZhYtzkcDeMsld
o0+mx0jkBw3zW03kxLd2q/8/VJu9CWCtz4ej0iIJWEHQiKysiP6rQhq4av9Mde34
1sNLfmAgl2VD83w6SQK2EyfKia0pPfAxcgKhS3JnLPxHO9Ft+nQDuyHZFuFMRHDM
0+WFAlG5s2ZeXcoOo2d9/8603uQg+C0UCZk61X57eeo4HDOva+dRfUGF1j93PtF0
6bfUmqArov8stRVKOqFFdsNDR2ABsz//M/yE2a/K9cpl/ns7UWPDgaG6eYayKFFQ
zGqJS8Lk1DDQTFz+jnqnoWm81NaLmUNRBmjq1HFrDXLLryptU4LLSfxYFrShyFdP
ncbwHHT65gGuvqeTEbBE/cf2n5WKObGQzYPJj3hRhh5QOOUgS9XCoH0Xc7EeDn3M
tGffkGvCJkwIbH1rpa7vI9wXEpnRiv8eqpr+iQXgV6mw70pnK8ql+/tTUlehfah8
FuE8jmc1whRzNkQDWmjluUEmhB9Lw4OtKLUpgm0gtWgZLbaEjRODaSzOoQpOssoh
p1pjh5OislndcCZFJXhyvlDdGf7idvHDr0wNt9dt3fIijJ/I/5xwuEDFl9PXo9bN
0HMEEhsW8/GNluVyQSusq4IHD00hkJ9NVcNjq2Su4J/mKJRLAIh/EPQTNaKlCccH
hQbda3vXrZHSXEd3bKHT9f0CW0ab80Ot37g+mN2mWaNvPMWM6xIM2lE645O8skIi
02sFG+9lMWqMfUieWPO/Ba9bT7Q3dXfT34q2MDLKp2k=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iHX7mcf3zDVp0px095DpihpONz+b0g8b7ZYd92v1Fj8OhLFi6Bmy8xEeGGlbj0Hl
7WJNpy4s5O+d7EBHpYy+5GIED51kZee56wl7ZmPQKm2Z7c1xErWOzniIc2W7OtDn
WcSIwXYyMjpCmKpBiAuAVMx85LHqHg8mXaUD1i7I7+a7f+kvdGUthVh1GrcPV1k3
Tmqu90ZpwF5rNoKG3i6PanZSRKfDwRHHMyBY5UEu1ds6DFV90T60Wf5OyqFMgiY+
uqFo40vmXR4IfmtEEnChEdYhbs1KnAL1Q4HO/Jv7BxV9f6s9Qvgx4SlPa+lEeVPn
RKI4IfglZ5KDlSCIWZnvCQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9504 )
`pragma protect data_block
Y+3Hg0EkhwZEHzNvqj3XD3DQLjxw4ekW06PJNy4Yp1IaTnQy/ScAhc+213SdVQE8
g3f6v1KZ/tj7mXTF6N2jGVAokI2cK/vAQN8w/HM4cgiXZ3EVxTgqvIP8kkYNxiOm
pfOqc5oL6IupVHdEbRIciueg6+djRjblcVXxVMqw1LBGFkW3P7XEna5e6c9ai7ce
tBzhudX8LM599TN/FccwCrPHAc4egKvOPU2dIpA9k24BARgM0Vhf5Y4ovhjyrhxk
TTdBZp6wGZ2AzAVwuFOYzrnr5PulsONzOPnUlGBS3KvMgB/FvBqvez4BEECSEeCK
SD/tRRA8wuEe2TkcWz3sjGG1qyTF9KmdYPiQucPlhnb+DKvTOZw2Mby/OUc07zhD
o0j0AiGNG5gnj+pDam8vTGYfJevnU22adt2NhmNMrx2Bx01QkN141oqasPtfiRTe
dfr3TTRKStcG7HGcgnb9x8v6I7X/Di3w6cd3f6ncP9GYNVbR8WnHCGH6opz4ZAx/
8aOG18wBN/Mam8PiWJdDV3J/7mj7qBxzMONqMNqNcqnRftXlBnpeznN3zvNiL6Kk
0fHPK//MEW+VBSDEAO0vsPgoRd7/X5OM+oc5UJQwQU+aRSSmzB9vUd9NwuL/InHj
mmY7n8ulX8YO14u+OSGQsO1wX3xa8jLRuJC4H7dOnftFBcWdo3wBjfl8Ha/oCf5P
BpScsGp4U27/1sxmxqeIzbDdUnUqOcrbvzv9qck/sphQ2bk3IJZJ63vuGVSzlk/1
SWsWbEd63KEpKiH+sVtcq3X1zL9TOz+3FRcTUrKlQS3y/95xSOMGAf1uwohr0an3
n54gx0hpFyzOHenEQJ+dISzbZtIJSoTQ5GMLJy/pbNgVXXDUo7ThyinubfZ0uKI4
8X5rBvB7p7neYraVwpuyR9DUu2rt3qO6o7GL3emo2hx06j4Kzc+3R5AXe51xtWmd
PMHQ1SU1TGs4PfwBMIisbnaaIg9jnAzjq+mRzUEd/2MIbkbAYjl0X5BCYMehug45
bB1hMYq1eUJmZQJWpoW8rn+GwU/iFjwR3xPIToHBzmLjadve8+CfPBaFPcPtUfnT
7DsldxIF4MCCKeZrY9REnfkbdEhbUNXmUAEahDUi9njsqtwOsp4COy8eDFEHmJj5
uROdGF5WHN6QQNJgRIf3UPLEubANowIg1b9iAgBYZwFK3FrNM4slpjEKQXIeiFdc
psPN8zzUoxniW260o2W/9vMpjFiOBXy9q7PYvYhkL5RyOhiUEsWI8efBU+MdFiqo
DFdJZQlDWcNrv4B0kVvLYPry+k1dsjRMn25LEVSUCDXs/2lWS1yd+yebsAiKYKwv
pGrMOl/AuzCk8C8VygJJIEhxGnbyGRtcPOpU8WXkbP3cH0uU8ooCnYc/NQGsbw6Y
WYyfG23RsZBnCI12WpNqkXpEO8oKWjuBAt1GqiKhl9vy7wInGUubep4PcFOPweYy
trZorDCMa1f1quVfj9XI+4Hys6yN7135dJTIxbhVC3fP2xlSm3HQLEemE5WWdR1p
FQNBTAHPxCyUanXO2C6u2+fmq43DHc25WnKXTByYxFT9vnc0oQdod6b5n+FXvz6w
VpBXJyt2LL1vrFLAPD8FKIXcSC1ID2LuufTEOpvDPtk7Ptvl6xPb2M8wrA5xGqCz
WlRnDGUaLUqX11zwMF7FjxFUZZcKbE1SbN3Z5Fghhpl5OEWwfkcVjbmDQJ23+FHb
5BsZNt5/xERqOwSp+j6r2bw0aCvFQOwf5DdwnjvVyFXvJLjX+tzhedySO+W4J+IG
QAQO+N/pyyPdmqZYCW3ry+nWki6ZKXzjy4HXysTlDaTrg6OAVQWE3esStwBRUb2J
1gH8qS7RyE/sFZS9TFLK9+4tHGSloGQ2S0aBixzD+Rluk3EKYwLvZ7ze+tIp7Lzj
4VbgIpOOODN75LR61Eey5cNk/t9VvZvBdObWTzRhBCtf96QCAEwWZkP/mGkvhZtV
jjJ3ERQApgYnUDtSjPBvuNWos2ZmD4gSS+0+wwAJ8lVejWsDdFdwDkGTR2s/HGiI
nfRZdgX8z5triajFesTAUG0xbufuCnMEuy2nHIwk9gK0WQo1XXu6CwqOwiH6EG0c
4RrubE2LrRpBFEIxr2DPrFKLyvi91p5mZob9JpepNIqQdIMQv1V0KIGLwXKz7q1k
K4amY/FukDGNIQ378Od5q3nihq7ijGWWtfdcN3e1qpjvXPYetzR5PTLtPSh+6smp
gZQdZl4pSf3gvR1+CREzijVXuTGO81KGSZ3EW0Quz9mT3vrcaYO6h69PhjhXYAJ+
No7tbKjuHAqfLiF8GoF+EnZUHaP/ypVc6ix5oN4dxw2HNsIKcaPnLQL+b2UIWSse
qZ+6kh9XjyhwSgeLoWelxOy7v3zlBk1SdZHU7Rwj8eZ95IdedPV5k/Ha2MOFX9e0
acbQnEXwD5Uw6uciuNEVdtvnQfuISYK7/mO9uWtriL/lN7vwQSoAaKWLbMJmKzX7
cpL/YPzOCpUISkM+MseexkQSjhmmY4Lc8qzYQj5aFJEbxbLSKxdfyqaN+b+ypD2i
Oo+E146nkeC/DeTDI7jr6hFx8PADXX3/16U9Xkf4uMJBRxYWmJMNiy9kdi0NcfSn
ntd2EeIkZAwVZ3LhPXtQWoaZSIHZPTLqRfcxc7vEcVDX44Dt86nfw+E3qfAr7nou
LaD+hmb5uqxXX4KsK1wkZa3RwNMNg8XeODL+f9SUDq6AWBKCSvqhPVHQiQ2IDf0m
vK4leZj6yikZdjvkab319nZsI+5eOGKGziSL18R1EhQ40QzNyECnkwrbVlMbvG9I
immwMXoO3L7UEP2pEqNYA9A48ptY6BIp1D7/3O52Xjb8/hel7EfxsxVOBv0RD0mX
qwAOs1emicaGqbHfhn7wQffk7SKgL+37wz74PaRGpKCntq9Ouqj4spfZrBy2uEXT
eZUpyqzps2Ovt+GF7CZTYYQoW2sNK+bdCBJtjbJW+8EW9mvbeGj/z8pXOQVm+xes
1lV3zgotQb/WJB1JOsaa/VrOE5JZ4SM0h/0Ki0Fj5FED8i7L8OvlyIqfLbtyzN7X
LcBcveeM4slYyKVfQutXGIrLpnl8Wgye0Rxl1OnvEp0GgQYMAQGb9f9gEf7bwL1T
ZCBICG6HUUNLjiZEYGlrCdTWxYelUwBIYh8qn7T0Rf32sTahCDHIN4CG+V3AFt/W
SWxmM2ZhEkQ0D6Jc08r20uPxtZ4ma3859v1cHxJWqiA4WVHlex5pUSrII6WNIyqq
qQsAUVenixtg6QUadJ99YOoFPPl0jGA12WRYadpuKk2+jj/F++pDIjx5UJp0MQmu
d7J6a8EvHLcj0Sojk9WD0FL/oiSK2r/jTJhaqwYLt+BFlF+Z8lrLPo/1eXuHYdwd
vzHhOM3bia8etZZ3rrnyVw+hyU5MgzDYMxe1FqLJn98rI+trGuqVCZDqPHnedHaT
cmZlyhp9GO51aSnwxmwsM+PZoVuUQSyO88ph2fvn38tw3g1mtLGyfXLRHs/dpERd
z/48XR4gyY3VQLRDNknRRXfJzzut1STjGWTuPgGQi0+JY/rmWEvK4o8Dw/ljYCGt
FPURVzzG6v+HQl6JgM4hv2Rn+UqbshsiRQN9zkamp2TkPfu7RMSI+CQG5YI/LNEZ
21/22dJavQUPsdGluFNNC79lKzNNrLkeBArVCjGs7lCUvHWZDwNS8QMMjPmhpF4i
jFfpLDvxskZojIN3eL7p/oSonfNQFKpZMbU/44PTN1/8PXoOPLBbJ/zcpaRUBulo
yZF7KD6TfLKF7oQRIFlKwl39do19tXfgqSzpO2zj5hNdfIY0yJk/Ck5NxZdPJTv5
kuB0ZpAt6R7nhM7+r9ObTu1aJBrcQvzThZIBHmWPxrmxAck3Itsvkgf05wwdKMee
aIh+a/lgLy8dVWiQSvn8fgawouCc864WmJoFOFYAsfpTyW3tGU/0mKpJ4eVAV+I8
ons5IRCHiOB58JKrL3mAvdz6JPPPLiz9MuIaTH4edTy1mhhLsQnMF9nyxdxTg9Ay
oNJYeuH1zp6CZBOcP8zhHj2I9kp0S7N+zYmNCtV8wL65cilZe12wpzudR7AEF1aD
kHXKpPIegamtFnFFry2R/hhLAo3ilMdN42tw4CzKEfL4Vr+0hA6mYyKm2omJCTgh
xfwaN0RHxWCZoA6/4GRHL+8QGEKVRXTDA6ElRIX3OzKxZxjisYLDExENUgFbFr5h
onpasuHBToVuuzxqoZhTPGupjJzJ26hqGSP/Mo/px5766NY0Do291tQ6o36+ISiw
lOQHU6TSWA4oMemmXz+HQxoiZapftDFjiRfwkNTl4y/943jFtZClqCK95O7gYpoL
l1d3R7tE+j2yZ9x0B9sD6G14TLQcaBq/ksWpJ/S8TCy/HTG2uplzZ+mZ8KEoxKAD
Bs3hPc3PZBodxcAbKVGUaxY6Vg4CoZFe8528XuMz2BmwRvnO9/XegtZeJ0ZjXidi
Y41jr8hcstOSJ3UOGcvgjjCvW7Dby1czcFs5a26jsYcTXso2ELbjlawnm0yjJ/d8
jPlShtkf9C3TIaKB7sKdVrl9O8a5G9pOtJGrHmYD7aJqW2yK2K5SqpwSvMtkgknY
Z/cMOnm1s0tolyCB3idvAgit/z0h3WfUEwTZf6DrIfpKgoeKy3R0Iss6c9iAv7u7
TCF8xXng2lVp0PNdjZHJNLU+8qr2ZWKeRp//e12xdtRt3P1Ih3Tk0tXdY3BeqKUo
2Q6BlKzXcmknR4ru/jgmCfgXg/+W8jcyOVNNmAgbWt3cES+OqdA0RUdR99ZuC9AE
OKaL226KfNozS8ComUxdcqNkYgvAinkPmzaEcUHw5OFonKwiUpHYtfrJu1I2wsUe
oQqwN3UTBQpMvd8zyCyq/16KWeSC9zQpSvpiE8IlBH6iMyZ9EbARKbHHIzwzMzNR
fea3S9AITFwddDgmHpEatgyH2xkFswqQ2vGjdPrMaA0zJfx1Giir25Wi5UwpeyRS
kHMXExL56GWapVUBVVaqzDGYyxnFaE6ynT1YvkUXt00okJQu0YZ1DoPaURQiJFUR
tHEV4+8FtfG8BLsfWn8ADRE0k0IJ5giYnNrEPecSJgwBOSWL1KVxC90DCh4g/bsR
5mGz0DTvfQdiB5cwOaSqjiA/TfmPzTBXrG3PIlAk5wiayqaa7M2y//PF446ikgb5
VJQl5cwNSSQb/Jxb7wFa4iDqBfvFCsXmercyHN1Ce7aY0RDD5r/G5hUGdM6qfiJZ
k5ivMNYP+rdDYhhlyhQITlUdbGifdWsulywB+lOacab8Ygo+C4wKd9YS76eaR/vn
JCgApze6V2VfdOCerN+y11lJMhXY9OaJLQhZWBs4uoqo4GUuXSvRUzfZJjwCqA8x
evmsqozim6Nfhg4IIBlgyvJdTATbJmz57BJD9KhFoC6JcRD+M18j26sAbbf1yEG7
SeCvyqnvidoEyN77QiRhf3P9Tvf4DlPA2043PEID+YVaYhLkDwnmooFUJYM3iMwL
tybfTJj8SJ80//y3dYBhsN57xzhfHyFEdXWkdSC3sYLlfK6YupLiy9O8Q5gzfZEG
OTop+bxaYbtMTeBitDa6kpNRDxHD8uiZioaDPLPNnsPNMfk6hHbDWZ04pahp+VZB
MJekWj2JLUuIslWNa1lGX1JOl/J4osgwBEoTcTTesFXYFAA4NJcxll7S8zfSxRTS
HmIFAKBRlvQ35QMJ+Tt9VeDXphxv0VY09zuEy5pUiy3H/Jtuwe9KCA80irmOF8Ze
GcEMKjt/QZIfz0UrmOngc+gupp9yX29ehN+BG5zQcTvJMXrxVTZH0c/kJCNWjYWv
EaCj4lJt4+7zpnMe7LGu+bxreXVLTjhEALxnfm3hZPsSeRuPoKk8QuH2SDN4dIuc
IbN6yjsOo5HcXM5a8cNw7LYEc6gxCoB5yJbpQjJzQFgBTiChe36g5XghJFwskPBC
/2IR0xwbWS3u2h7RyMQrVHxFUQF6jDNFMMRVde+Xz0ntsk6g73Y0veen3VigJRfK
VX4cWGgQG7Hg507yIWZYQR5UdblMyUo6pOtan3+3QqruxUd1nKvZ+zvixec6u0BB
7O+aG8UjMFNj+na+yXOP+dz39NGJyA/GbwOhde4Oy1K/VrkhcJazbL//AUGWOgHZ
Y5XqDxK5i2P3OOCPk9nuadp5kSacPFa3SHH1SUV11ocukq+03LjSIT3xkXJOkWFF
lnnM+wC87/mR9lvrZu9eBAEhNInQBtA/xh8y+D7SMHZ3Usc6Ay4+74o9BtUKQ8S+
TzEmT0txiMfgORxIsnJ1/zpk2eUFarfjwY76brmiyH8hVUXxCQdSPkQZnZoetjUJ
cVGlXKOWwaTKcg59v9xq4vxsY7fVqTqISEdx1FRKGXujaJScW6KMgIxBjiSRWvTQ
lromLyW6X0N+WghlQikpmYAt1KiPCjQI8KbGn/DN0FIs5/foscXjE4kEalv0A/6/
ZZfD9F0oCuI8GeFGEGQzpMYzZhzfbDj0kVurR/4py7vJwbG2H0rtir/fkh9FOl9j
z5bvY6atZjQ3m6+/xs1ly30FjvXWjz3qCt+XwTfuSZNgvYiO4pWCJZv1E005ofwq
/fWLEZmnD057u7iQysSq4sY8Bu7wlvbmhZssiCqUuN8Ss3a2o1Uxh7759kEgAKKZ
IC77RD4qgG5cZn/hj9VRpfNGmFgvTKOi6zeP/KPu4fzSQOY4949u8ghBRMnOJvXI
AFAMerJAhu1/6RehMabgIxfvJZ6ua/o65u1Z1GlpA9ZK4lll520E6ZahDLObIwZf
TNDeohxkMOk6PbUInG3sHJkW4iYJPq0AGEt1VOt2EGR3KhNzaSKAHu+YXJymvMKg
NwjbxImQfXQhDxpn7jnpSLrAM26lYFp0ZMTmXW4paZFHJ7FUWYC2Z+aCoS/tdvMV
FLyAmKyJSgtvkkTbh0V3poiR7JiN+CAAf+qVuyEmHVbT/J4xWmZPVONMNJBAfwUt
isIk10OUkAPDZ6jUsvDi9f+qr7XrEDrd7t/5AQgDKhIVoXUWakmn1gq2CahKMb/8
guQYmZqOytz7RaRdK4Jl1J9jTxeJ67XaEwLCdfR2DfhpBNrYBjoOLj0BNRQBCqWO
UrJREcAv7j3/5sZu+kLlKdZRe0SB5JXwNEW/5ZEESv1kVNZa+ubeLpF1mNOYgFa5
03+PdsPYPb7cGBPcGz5w9dFm1HSUk+7aHUfZOg5fIWPe9EkfrWCk4HDx5d3XAvKu
F7vtEIDRRBT0rb+OtXWCe8Fbc6usTtsPcM3Tf8BtNhvkvQJBbzkictAjUygBUSVN
nx8olN4JXmzIsXRYuvYz9AI7RihtChzUM5e/f7GrBQfeuL9EBexj0qyLRUbaAQ6H
HLHNxc5YEKyR4yRgVdNAx+SpcQHG3aqo89nWaNbfFoTNfP3iUCZvjvx8rgUUVK4E
iJG1wakvZo6TXLzLp5DfxiRiZGhnZ5vuKw2fP0b2Sm+EkeThpaL9ytewreRDdjAY
h9lRGDJ6DJYu4jssxavdOC/nv5guJPVurYzt742YBIXuqUsa/9RKxK9e9Tn8hpp0
O6C0XoEhMJu8VRYqRDSsRhqAJAI4h9N6pP2RkTy59fpExCUIQAqbdsGOAMfOCg1H
6vqKB2T4nzPTPGpQbYvUqid7ONfFWBxyU6SJAwuwvOpQFNL/xxX7OXhWB17WgCPF
ULcxBt7wTrV36gtquYU6D1BtmGw4dpJEoCE/BIzcOFkMlaldcwMSraKs2ew0E0ig
WfXxHZEv94cprwieaQWH7aFcU63uzKnEX5zUbwlUwvtkoUzWojiWWWe+AfHhUfBF
KQKVd3cxR8NYxL+LeiFshY+9aZ88atFBJhHiq1R82McrYLn+0SXN9GvoeJFKAZs4
Bm9RUNGjbO4cxhYViC4kWdNpT29VMITbfReruTSu6117u7byprQh8sAw4qdVnqxF
kWqg4yPCcSpfO2fpyAKQ9wjdbQ3Akw5oIzMGfXYKKOmq8kdayjQfR7sLY3zfcTuq
yCQsjxFtQWYy7eg7l4i6Fk9HvdG4GmW6BquNO705mqiPh2bb2q0CNYesCJuFSIvq
Q8wtuzAXzVhzWG/2JBFv9JA9Xo22kZrMd5i4jP1+cT+CfHpYkgBkE2viHZqiiFJZ
wyDo7ey8e44f+88SQeyEv8zT5w0yt+1+z6NdpOlQIsCKuueUzMR/z+mAsERBtiHU
oHW6GJrw4aFCRHU7l379pwFIaS7riu7LJcnMEH0GPqu6nVDGC7ZgeZtkSaQjAY2x
hyZGi7W2tN6gRv6Wst0HGSfIZp1xkgnWxoM5BQQG3FUGvxnMFqUFzT/etwiP8u+Y
brHzblbwrbt5pKPVQO16ImxqcpDsqL8giB/4yV2wM1qemmgfMdDm3Y6MVLm9CRwh
Eeps4C5sNz9NPtMW9bMUMPCoMk4ki5TTk3kCsUVtRiwdCJ+EsHImWTODgEryI+9D
VX0RJ0Svoya/Ir9dd7btYKNXAgzj5c3ANP7Xk0tk5+Auydxe/xcTFPk3THQVlG9C
AmEof9PkP6dsbb04oge9QQFsa7siDdPDzc158gA5zuzA7XpHRVUhqoQFuzcKCznT
j98DFuyCEPpWS27z9L27epuEjUGNUI3dpha3x0WP3T04ut8BrvCBQrEI1QnFbItu
r635a9Kw2lRi72+BUuTtC+G/+neBaFWavUatcmUxinFX0YdCdp+oBLCMlQ4pgOmY
oplGu3QfsrNLlEsZXWhRX5tmLR0RnpuCejZyihEgatVm8iw+G1vF/1+hm9OPrZzk
767LxHiBaK+ianQeMtvutoeD1VXop+7rc7anvatSpF5JTGHUWO1LVyT/ECZgWO4L
5IUZ4bQtpttSipyl3IlyTF5jC2WYperBUMQtaU8nYUsWpJ7N0t88Cb1yuacNpZ5g
1YrRdH+84MBqJ48x2F8mVH8drD2O8bHL/pfu3IV+dxQIBbq+T/R5xLcgl+KqdPC8
UmFwF2CjN1QBVpmWn6bkEAfqLd3RvhkbA4z+691X8ok5YaW2XlYVG4jG0SlrZj+j
Wi6TFTSh8qbQx4ZnvAhFHieCxp2HjgkMC8U8n17/f0+z8xt9Mc2hUoUvX/ndq3uc
9k6In15T7tAZuBTJeGvveqq9nV7v2KdLtzKI0WZqFWkBYDm7H+vMJU6bXXh+FUsi
Ap/oqrGlcy4Gsr2JEwpCR5VwCm0JxDVdDBcjxJMDKIzY8RhmLg6+8sY9pJsUFFqx
YX133SkJ3yO6Fq489wpTXKResd8q9m7mYuVn/X+55oBIna2ERDD43xan/RbBKYnl
vlt6+lMR1dD4YRncr/SrZUDI3+mPS27ftgoj4ogZIEkdXZOP7VfdoBhq1vlR9uMh
KP2Xb4avixfF+29EvQRQjT0VjCqb3Rv1Pm4cR6M2p3UnKiDB8Bw+cNpLpwnujXfH
YKjNGb0ufIPmtJg6G7jSPVDDyTj+r9nBeOijW1+gMa5pFJ9TUEIf95VAe1cnSxhj
LiLmVxgH1Y0EKzzG2mcYa+911mmS8JFLvbGrfBW4V5HxayDCWIjyLUE6oY7eRz4U
940bvFUsvqI8CkuMJI3pSgH2KO2zkmwWK3MwBauCR7UDLixwVI3SGdDx425TaoQr
v1c5wpbCsXT6aVSF7fsicjT3mqZTJ8bAPQzLnR2mtqk3634EfHhDpDZ1w+obIXGd
Kn4qQDXM9RR67yxy3bFxOwLwZAwL/Lf6SxSepQS+y48bs6HrNjMFXMAx1ucvwNcF
uIx4DBJOTyf4THoNWHpYUmfHbVI90y4lZjYR7sw0p/K3ZrtkNbSb6YZ2P1Fyj2Gv
Z+wR/d4KS9BTXZ/JzKYLq9psGfNUpqVHdVZjw+djb1gvglhMSUSkO5qXBC12Xj0l
vPch24zyZTJJHLyykn6y76w4gC+rSy68OpvRtV3lb1JWjdsQ4jr+L7Qe1xHPIKZB
mFM5zOn7SfMLJ9H3if36LsgJsPjpKmdMvieqFeK6+CsgGuCliXe04ztiV1WA7NnS
kZImDvJBMPnX3R1Gt3OemjIOEyC7yMnvul5t9VIJn2RNYEcFZ8Ssjvfw0lWAEP0+
fSVUn6fIaJq4lt9dguaofhMwJfOn7WPTCgdE2vTcuJdImknbQot7S5KjmTkR7TuW
0o9Wqo3ywhLONgXPRXs2iqlqeHGflGUjRpL/bpJQ7rXicDzCZ0EjNv4I/1DdfVvJ
tLf8r7YcsDpwJpVh4hk5uNKfI1adOPzPqNN8VeJB/R26+IWnahOme86hOMU7qvdg
ey59fsXWd08yRcszO1GMl8ER/5oYWBD2/BCDqvAVpQcaxfFqLbriiyBX/8crInqT
Y/nTiPd0u7S8hou+pjx3Ewjq2MQI3GPr5HtqvyEDSyZkvP6ZX8pfEbXBkfPCeVrE
N4sHlP69roBV1S3gHcyv00T04EGlprQdbjGvrzmfRYoyptELiW/OMPfYEKkcrn/o
lrn4yvqVEJYDpRLMqa/+/bldWL/lFmd19VZf60HwOhobQQGpBhxZOU/f54fqoXnv
TvTXI14vCXy4S+Rs9cUBjTAkDOvCb/4+/wLGBGfL+oBQ4g22nwTxHS4GxaLsCsFw
ab+Q4iMqrVmGVN9AnsZIXDtS/20QpCGILvWpm1j8WEUlM7CvFAi89sEuztnRcLz2
0jHtXBP/sZW07pAY5n3hn1uP6G8YgjUQwodN2ZZSjbZs2ZatuBryMWqwKRaAOlHi
7ZOSZh0wihr1QS9/c94hBL1nxZzjoP/pnWDcokelN8s7fekAOu3icrdb6IQR/5Jk
30kLKcQMsghadtEIQHe/7UbI3oBwUq0RdOuoeGLubhU1sQcZYx/RyT7Q+mdIJzM+
rj7euAD2T6yDomH2ht6UzKwPUjJM1YdyGad3Qu8GRSYMWpVZW9xm1S3rMUMyUi1n
dqdLuV6kemuWu6XlKvsQwxhu/SotTrOKPrA0aXrxzplq0RO96omdwOesz6RTea1o
1WtC8JwIsv2mzlPw6nBLupPd7xlxUES/Hwq4cYhjnF1tbDNrCtwwdnzrtQM+hNIv
1WLzDaA8kHkpdEQOEaRmMPlq7EnLq6CWS4EfTqCFqjHjQNn5uVSTDpUt1gU6rWH9
5WxK21Fd9zpaCxptr5gBzjse7x5UG1ZyYTIvrl71DCf1xBGKiYEsAAvKqF5ZJ/WY
fFmlbbFfLVKwYfu2WJAOSC8s4twldPAV3eGshI7y2IzUQUGgG9NnZ6/BOobBSfjn
xLsorxjeqi+sEIwm1kC5Gh6CaOy+rJt+uJWSfFShcURtcH7OQ9dlNV30P6NmwhxA
bGMln6GdzPJoVIw5/RZ37f6g3VDB90WWrbnsoDxZxUZSL5nTjYcEgsVDk7QQwHdx
p3M3ASbdqmm3b+UN1imHaAOp8TexAnmUt0HQmbaR44FAJrOU0R/WaZsoqAO4JDwz
KZOiqaIiXHmL2Kj4lu51DGe0q00uKlcsMQgpY8UIxsFGCaJieZjP4NkqZoYB7VWB
be3qAEBhXTOiqhWS6QYN4BISlmTe3GwBtBjS7sJh37AKdZboXkfi3BfT5h3SayOP
B484U2JcEBIMhRnUCZzJ9tiCuVxbdsm3p3Fkj2F6bnJpBNfxHEQ5P9MzKQmbT4FA
uMAqTkBieGOAOIVzLn4s30CjzW+qrCav4uWTi70gaY4AZWkvFU1y0A7IFT63SUn+
VzUie6hlEhiho7e71qQc09W7IcXIGsvVORx5HK9UJCtLUcASDssGIop4xALoRzfp
K1YtzFa0ajoLrTQp+X/rFiWgwgpya3+wfDWl6smw9ToGm83KbdH8xNN/e1/o8qx7
nsOLIfcB67gzlicO9sZNOdHuJ4/HWIvmO7pIM8RMBQnDEqUJA59Fl4GGuRPg2V2V
isgWIOYkOXcMhjbf0U54riSul2TVH7AHQ5sfuUmGY3+UdDKQfI648c6HJHE+HJw+
gT8ZME2xmkDpCwlcn10+ZmCnApEPq9XVYTBSo1n3JDyS2d/oNK6tzA9ACxnDhMH6
KWgMPPDvRMh+ZstwZj6YBvlGrgoTOUiCy/8jpifoTjLl4VjXnS3lDwM4UCyYGnW5
EFwTs8EWpCqP+Q8HvyinN64+1FNSwvlj22UJPCWBnNlsq4oDQQnPo+BClXJGC2My
wHffi/Mux3LNJtoh8klxXZLHQ/f0HoMaJXIkKC0g8JYvMwkJNp7YuAId7DApH3tm
Yt5i6Ty3ecQYn8hcdcX59W/9FJG80/2HgalG+7w8phMieMJcGOKu+AOWyrscyBvf
hRkB0AG3wj6rkLkbdonoctteuXWYoLDCtE5hEZkXYP37Jobr+cSj2NdVvbMrNQtb
a9PZoL7MM2F9xxwsQ4KNh19DHKI7EL2Xj15mXhk55V3f++ZlcTyB/Ro68c+Br4R0
qusujDyIU+rtbW++Vug2ZwK70TQsqNRESi/glpI3JQrfHWgLNL/GH89cqyxXR98v
JdtrAsnwWxgjpj23+kBI4g26P/d3kC/XRuqYbQqhExMWw/pawzt10H6wwUpcWLzX
bU5roI1EXWktTl6po/T8JQal0G1Gfv+P+g4zb4QRiRwoP8Y42/QKi3F6JoaK8jqv
0vdHnKTD/1betFeTGeypcMJNQvsxQv9jjD8ak2RXmn0FxnG1ha3sLo+QyEWP4AH6
O1mYhyeRY9OK7z5u0Jmja3o1x8ha0z5GthQ90Hv8ASm4SdEexw6bOd7IK8fPyMGj
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
f8eq/uPKF9/r7PI7Eb8xvrL1TuDsTUThMfYR+pgw0lB1LfLvRjUlkcTmh3FKpkF6
f0FNXltS/VtUbYPwp+nVlFVzcsbBNn1Fk/fqrY6sQd7HAE+Wp6Dd2+TC5cYqNWgL
cJn8hy1FJpLziGBbBbY+PknA70iu+++2089HLmL2s+5HOqbCdbXE0xfYEaJ/3PEv
k6aMaU8s0LUXqet6pg5Ke3Xo8xI2K56bxNCeC3Z8mkf0xLcR21cep0DBm2DAzShi
7YTLouKQo5z/qhPz6GCqYxOjKPknTSWGvsrlo9qa2bOrenOgrxM8rJhsOr2DXbKH
+iIgcWegoHcLX2IwcwpkUQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 944 )
`pragma protect data_block
9/WfDK5gQ0tqrl8+aBHsNuHee1UVym37mfs4mRBuqQsBO5I9h0kHxvhYIHlDwAij
AphauEj61tZWVjc6fTWtuiEz4mFloIP1mZIuQUZplFdTaUh1hNvy3UUcXU8UxTK6
Be5vtHGLf8MDh09dkmpoW3pLvdkVAtTVjjjLYJUhq10OaiZ/Hgp1i951VikdE1Vs
Z6uA8vQU5e46c0ZXn21ukVCC9EeUcYO1b4///XOqJDM8jrb0pFtL+SHyxt2aGY7c
7lJD8Gk8Q8XpOIt3bmPdhO35aHeHah5nLngnDrkn40DBjOPpR7DoCRdHe21lNX42
MGyJxiFrb2nnAgjn+BIZ/CnsPjI9sLJ3zfNJEOOPoZt9A47xLjmdhJVI3N7Vv9qr
G9tfYFCgbOZrRk4GJDM0Eh2Zv/em8R1T75MLG7bSay6BKFQTVrYYKIuHex48aQTn
H3L0tpX51qjLfshlHwbxsLAyshzDPw3ibM5DwDQAfkyvv+IenritJobWiVZifV5s
1EDSrsNO+ELRwZGPNw916Tbl20uWszozR2JG6KHGJNNz4DrPyalN7cqCoT5hQWEJ
xC7fejEMaszCD1LcAJr7v3kqRz8sG+aqiHPgVYM5ts8mz9BDwL5ptVXbLJBwn3+i
L6hEEoo1QcbxcJX1Utt6g5Za98xBU49R6QvU6aqwWUJXjxid4SyCTUalThLuVHVz
9T+1JmExdxwofqFadAQgs+PqBz8DLQDkhBikozigef5xZnieZHY4Ec/M+C01b5W1
nwzizQhXt/r9+JmBHjRaSq8QqkPfroPdyxOepisuFhAPbdMcfgH4hyTrwE+aMZUL
4GJeP9hKl5c9G6EpHxGpCmBGvkbCu98JtA9hepZN8RnEbdhcEqpQEiZ8xG5vz7An
g3heLRg2Xzg/spbsxVhWVwddgVHGvH316savtlCbcZWRvfwlmp+Cst120s+xbgTH
5tAYjDe7Ybp28yVxbHixD0EvnV9HQ6bxbufcCsxA4YwBm6LdVpwJuEC/uRMcCb+C
MEdcNmSbV0QR0LIlyhUzto5ysmEiw+Ten+iL80EIqhtfBd5UCongg985aktcBQNq
s6HoOSe03qh04NqLRczHd0EIaS9oqbyyyTde6G/m4JqTLlfFqk8I8nSK57oK6ke/
jNqtbpid+6OX+feljyk8jFfrXMaByNHVo2iuovdq8Hn4KD7FJoJ7RMYpeEbybvBf
T24B2LLeMKhN0fhTMlfU/F4+ffsI4hk9dtFBiVSjiR4=
`pragma protect end_protected

//pragma protect end
`undef IP_UUID
`undef IP_NAME_CONCAT
`undef IP_MODULE_NAME
