//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2025 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = csi_rx
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Thu Jun  5 09:45:38 2025
// ***************************************************************************************

`define IP_UUID _csi2rx250605
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)
`timescale 1 ns / 1 ps
module csi_rx #(
    parameter tLPX_NS = 50,
    parameter tINIT_NS = 100000,
    parameter tCLK_TERM_EN_NS = 38,
    parameter tD_TERM_EN_NS = 35,
    parameter tHS_SETTLE_NS = 85,
    parameter tHS_PREPARE_ZERO_NS = 145,
    parameter NUM_DATA_LANE = 4,
    parameter HS_BYTECLK_MHZ = 187,
    parameter CLOCK_FREQ_MHZ = 100,
    parameter DPHY_CLOCK_MODE = "Continuous",  
    parameter PIXEL_FIFO_DEPTH = 1024,
    parameter AREGISTER = 8,
    parameter ENABLE_USER_DESKEWCAL = 0,
    parameter ENABLE_VCX = 0,
    parameter FRAME_MODE = "GENERIC",    
    parameter ASYNC_STAGE = 2,
    parameter PACK_TYPE = 4'b1111
)(
    input logic           reset_n,
    input logic           clk,				
    input logic           reset_byte_HS_n,
    input logic           clk_byte_HS,
    input logic           reset_pixel_n,
    input logic           clk_pixel,
    input logic           Rx_LP_CLK_P,
	input logic           Rx_LP_CLK_N,
    output logic          Rx_HS_enable_C,
	output logic          LVDS_termen_C,
    input logic  [NUM_DATA_LANE-1:0]      Rx_LP_D_P,
	input logic  [NUM_DATA_LANE-1:0]      Rx_LP_D_N,
    input logic  [7:0]                    Rx_HS_D_0,
    input logic  [7:0]                    Rx_HS_D_1,
    input logic  [7:0]                    Rx_HS_D_2,
    input logic  [7:0]                    Rx_HS_D_3,
    input logic  [7:0]                    Rx_HS_D_4,
    input logic  [7:0]                    Rx_HS_D_5,
    input logic  [7:0]                    Rx_HS_D_6,
    input logic  [7:0]                    Rx_HS_D_7,
    output logic [NUM_DATA_LANE-1:0]      Rx_HS_enable_D,
	output logic [NUM_DATA_LANE-1:0]      LVDS_termen_D,
	output logic [NUM_DATA_LANE-1:0]      fifo_rd_enable,
	input  logic [NUM_DATA_LANE-1:0]      fifo_rd_empty,
    output logic [NUM_DATA_LANE-1:0]      DLY_enable_D,
	output logic [NUM_DATA_LANE-1:0]      DLY_inc_D,
	input  logic [NUM_DATA_LANE-1:0]      u_dly_enable_D, 
	input  logic [NUM_DATA_LANE-1:0]      u_dly_inc_D, 
    input                 axi_clk,
    input                 axi_reset_n,
    input          [5:0]  axi_awaddr,
    input                 axi_awvalid,
    output logic          axi_awready,
    input          [31:0] axi_wdata,
    input                 axi_wvalid,
    output logic          axi_wready,
    output logic          axi_bvalid,
    input                 axi_bready,
    input          [5:0]  axi_araddr,
    input                 axi_arvalid,
    output logic          axi_arready,
    output logic   [31:0] axi_rdata,
    output logic          axi_rvalid,
    input                 axi_rready,
    output logic          hsync_vc0,
    output logic          hsync_vc1,
    output logic          hsync_vc2,
    output logic          hsync_vc3,
    output logic          vsync_vc0,
    output logic          vsync_vc1,
    output logic          vsync_vc2,
    output logic          vsync_vc3,
    output logic          hsync_vc4,
    output logic          hsync_vc5,
    output logic          hsync_vc6,
    output logic          hsync_vc7,
    output logic          hsync_vc8,
    output logic          hsync_vc9,
    output logic          hsync_vc10,
    output logic          hsync_vc11,
    output logic          hsync_vc12,
    output logic          hsync_vc13,
    output logic          hsync_vc14,
    output logic          hsync_vc15,
    output logic          vsync_vc4,
    output logic          vsync_vc5,
    output logic          vsync_vc6,
    output logic          vsync_vc7,
    output logic          vsync_vc8,
    output logic          vsync_vc9,
    output logic          vsync_vc10,
    output logic          vsync_vc11,
    output logic          vsync_vc12,
    output logic          vsync_vc13,
    output logic          vsync_vc14,
    output logic          vsync_vc15,
    output logic [1:0]    vc,
    output logic [1:0]    vcx,
    output logic [15:0]   word_count,
    output logic [15:0]   shortpkt_data_field,
    output logic [5:0]    datatype,
    output logic [3:0]    pixel_per_clk,
    output logic [63:0]   pixel_data,
    output logic          pixel_data_valid,
`ifdef MIPI_CSI2_RX_DEBUG
    input  logic [31:0]   mipi_debug_in,
    output logic [31:0]   mipi_debug_out,
`endif
`ifdef MIPI_CSI2_RX_PIXEL_SIDEBAND
    output logic [15:0]   pixel_line_num,
    output logic [15:0]   pixel_frame_num,
    output logic [5:0]    pixel_datatype,
    output logic [15:0]   pixel_wordcount,
    output logic [1:0]    pixel_vc,
    output logic [1:0]    pixel_vcx,
`endif
    output logic          irq
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jSql9oXhGM5BoAdsVdGWUKacbt1IkaDcQPDllL6ZWQAaGZIZvQToLTC8BEwcEcPu
O84wWmz3XxicAeqxhNRDp+zZsT8cABzKrNcMAmqRwZMdmn2YMFMa03W1dlI0j69v
5UgsB+vIcTkbmEUMvVHu9C2SWO/7mMG7U+e4UBJ6MqSz+d8kh/QDma6Q7Djt6bn1
KNKN6cBQrryQM6OGJehNBJH3VKn60KfkfWSu8rF+Rs95yqsRE32jZy7eYblSdKFs
ovUz5kCAPbkN8vD93JklHYdWZRzbzHWhc/cyd8er2pr+osbYTWn0+2f2/SXeybFZ
63rcYThmcMYcggtQykVVFA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8896 )
`pragma protect data_block
jad2rPEAULlp+AyhRgTqHs4kbISOe5Bd0c8igioLhY8NjZhjhhh+d71qOWANddvm
wuT+DG06P88VlfA9bpQxJ+unjnd9fYbAraOO9mpR3hheR8+Wl/O6X09a/CXJYM2N
YW17YRYyJ5fRbMSHDwKKNaB7ElUcUvCtYsnUH4giOegicmUFybyORvanrAhv/Y59
Hrc8qAbehiLxZDnflOKV/ScXAWAXCEj4YAmWIbQvDVFBX/rKxXSGEIsgqmsM8aAQ
4hRoVcZXMy4/7YfRL5Urp14vWpqrIaCO48iaM2IQYsuhdBiqcq6UOYoQmmCD2iXF
K5VI3/NMQ/uSPPqRO1jpxhJQG2BNnn5EahV4aFliTYtZ2LkPjnuOzyZD1KvA+GKN
GESTOuP6AmH4Xu9pnFGZUkk38p5053LvvmfFS5QlADYurjhE7CQBeaTebtERYG2j
QtR4h3b4e6icnSHyDkTCV90ApGF5gaM+AbcaIb3hvg8qPvuA4v2LliJWkQTDc4Up
lGSpo0ZNynLgyhIBmnVBqfzpceCB56FLlY3RNa3F0iYEwhDuXsT8Z0/vtkLaBLA9
fxmvJ8Hq4okbiPvQTaCpdZ3zaWfrrwRCSHo0GwVBXB6EAKYOXI6IMTAVCKUrfYQj
ReqNg3+/sMxUDkr9w/HsI+8gpXTJuyktv7xIUYujbPKE8gVLs3QqUK/SjuygC4m9
VU+GqSvOeK+bpxVZTIQNpxfuhE6OjLiX2fecLMgyv7C/XnwfGcBsuJ8IxxKe31b5
0rv2RQiwUag5SAVpGLjfmlY40X0+Mrt7h5LNKLG1QfgayjZV4xFqNR6iBqTRGnyy
fqRHg+m6nDnCxdpGUUXUkFGVLcevppDiqMf2/iucn/hLuGPRmRUUO94IibzBsZcK
gloFhc7Dlab4N83L6B8N23IDAIu4cft60pV950iZV1bJFjtjj2gXeiM6Obd4NnRB
Vi5n1d+M35/luDMj3MplP9qS3Z8bvEef7CjgQp6EtR8l0adSc2cRZrIoM8fp1wUK
EJhxovBTwUUPc6q88wppqattxne5Tz7n/YFMdm6sI+UzJu3S4hgzDiQrK+Wv8ZoX
dXBvoXHJHR8bOHwW0M1Gh+hc4/XG6oaX+ENNYKfRSbCx12EWhrOhNKADQHuTTeJG
hVfS1QF6MrI18ZcH4n37PoNgYBuq7654sDQi/mS3ioCQHp/WUzRRImbHst3ZVmpP
UcPGgjKuz7SYXLuXF1W3x1f/HHhUomPYGiKAYDY0/EizdqbUnn0CJPxGplUHigWf
kr4p3Y4AoA6JCZ8StZTvrLFLARp8U5M7oG6vpwxtue/XwtrBkJd/XYb2gluv7GJ3
0PqIvqScwlXf8bDfTAsBwB8II4L3llbw9cp2Rpit51GC078OrqdeUE87DOlCsRX9
UJX/z8orSaabkZ2bLSeekM8ynRpZ03kj3Y1OVUU+8InR42V4ZCi7bH2LCkOe9iws
IQJ3Tcv9qJr6KGirC1WfCGCHUZ3fi7atKVlhxfI3XBY84PFXOm8LU6nTTFwSh6o3
Oj8KYKedV1zqqU7z8tXumxsG8XhqnfJ+HbcAmujDq2cDRYaNBaLWCGttr46vHUs1
JSTFwc17rbyGiCW4/Xj/i+hIMhywIC6tvYLAgK+27Q4wSFweeyhwRgJj5hLaYgqZ
J6faoE4/zqovi49AK1d5Fz3r0iZwa0E+t79rQOx4tGchMpnzEZSey35li6Bg2RAP
hWL1GYBIcNVJPrzXLm52CcH8Y1KXoHmFYusP/9i8BHP8VpY2Pg0ndPHMwuAyUYd0
6mmvwR3AiBjNSXaXcM8QcD4K1/fHzPXZlQpAIFUNUxZF8ICmqbnfvqPCqTco8yNx
9s2zG0nog7v85lZBpPobnx6BUtwfyE0RKtP4MkW3iT+rzYOmpJUODKf8iI0K17YW
U4+q9HmpNlZXaDEPJw5HAbrLg3crPw9xRx6fUcpPUJt/qK+N7FTIQG3k3PcQMHn+
AZt88Xhz+zszUnuiXuKhPITNwNlrKfPd1exDPjwf303JVIf0O7snadb3yvMVowat
IA9lI6KNb7eIHsOITIyPx4xMh6NnKdY6HCDzcWNV8d0XAUul1j4SK9TAxQD0tYQk
B+if+iA/xhHksvxyaSEcxHoOSnl9Ls4w4+r0DbCg9NFJztJkNBDk5T9s5RJm7N+X
Kgv/pb5f25gcbOoUBmheMsxkIKA1eN/2dW3xmXWP0tj2Mmq5yQOrn8ZSGUPB3bYO
sKG0GXdWOVKTO+PRwSfk3p0tOFrciHK21dTsFzzD4GqHIECNt45jr2/nQu8P9ZoQ
ylAxzjURBEubOhmONysimLDqO65qce1qJdE39mHuRX7ZmXK8nM8+TcMkGSmDgBqf
z/49vMZowft6W1lAyZmbIl1ag11UKn3H7kdnPgS1O93AQVlF/F3fk0JsaSEs1Eim
mJLAlLw7KW2yLpQP2272gdRC+/UsWmj4XAWiq/LNw/ZU88iBtrFD7tTdLy38QevN
lO5FT7sZY5TuLBMfjUPCChisxZrkqOY+2pi1MaPMQpRbXSND18a4/ohpUDBtVz/a
uTYcAITPQ0x5kGeCyPlhUY0L88egDFcF1dM6WG807S51FyJh9N5ifKZVMybqsPrR
hNo2Q/lqMcAVJai3fMH0Njl6jHrWmywQRFn5UxPJIZ7GJMEHMSxChMKSejp9ReU0
GaM/pIsNAFptZAsAQ7VsEP8S8f2wG94EqVU6A2alcCuA02A06qEY+3rSuzM7LU87
fdC2P4lTLauyJ6h5u2f5/iK1oisQvAMaxs3wIC+kANx3zni1swGHwMX2ocBviZfG
NtIoxT2kIw79XdweBSYQOftE9nZnNvMAZZFgZBXTkwhjkwfD6gd/FgWsReWNQPRZ
r5XaKPXaRvlIILSQAFqq5NLYSzBTTPmnJvLpcx8ir+rYrG3mndq2OGhByjQaUt3E
G4YM0LuQC9LjRgkiqrCeVEs5bdC5dSF4NPTxuZnfDOOTkZZuf6W+RqMfOgmRJhx0
YOsfmvMKJihV2c9ul8hmQHBvlIcjuYXrdco9mKWaNnovk14B8s4wkMyiWXl8k+I0
v1YBLW6kMUmfPZHl39jIWWNexYeJnacv0fXderz3ciP7BcLRAhbqHhM1yjA3Jk6I
TM0WEFzpN3Pz8dCK7T+ADcqH725xxY2bZRmNCyKEGqn0fYp2OIAfVcfindiMkWf9
2bo3O8pUjfik1yJldfARtWZe5ylbsG/piYyBXFvMxsOF4gl4VBEhGJH6c7igUvu+
avUvnjUesxADTHsVxkQPvSu6dxD4Qo6cK4VBEXl0h37ey61OKEXH/OaWNiIgopLq
9iKGgRlJ561A9Oiz62ehLcu27MygbsCmBRTdPifpRQviJDkITQK2MmM20YGROv5M
ch1Sog9Y4ZlLWekNNz/qAzZWlLVMfbNPndFKt7Lv+YySi9POIMDRWzDoXOpRPORR
CzYS+1H9goB/lg13NmTjzoOwDYn0/P5mLmjcmah0xhegYixqWZxUik4JvZQVrOqb
MgUz3IliFHzFWfVNGyuOsqH159QRLVo3+KLk4HKODHr1RnJorw25KgHf6GO7HVPF
1g47Bbr0IeK/UDmwIBW6ChtBwraUSklSbVJ/1L7FJAzshFVDZEJt5ckfITzE9I7s
4LycdI2Vkkb4jOzkGxhT1pnp9U1OcKI2dRKFb7N3m/0+L5uqvi5TDI7Wl8sb+CL3
eC7pqoexVM6Bd82oLPLzosNL7uUxIm3Xc5EULjz4oA+NPSd6y+sS097nzuB7xZ/E
+IDzSpewo0ezySmFKfPe/vPDsmmhW/EU4Qxt4JYmunqDFXh0rPozTqhqIYAvp8wy
HZzSF2T3D9KRJGaKEr9Ea21P1QtNTqmFG/R2U8+62ibrNpE4rDWDatEYpBNWQp+z
R6MHTtqI+MK9P4GnNlS7LCWnzok1O09vUOE9Tan7GlWlVJuZ0UhkIZF+YsWKVc5W
wOaYYptgAU7iibtEbwAxdc0NivIbrBopk8BmufwVRPxccTowaDACYBAtgHA8B/6v
1WYpuqdrnVt5meJaQ+kTN/GSPx/6IssMGyV4OeApt1qPr8ZdiorkVVXJnkFTH9E/
HaVl+FGgWzTHMXfF/UC9dowBjSOHqJdBMEn5NDdsUIdlFWAJQiciTsir5f8Kdbiq
XXmBYcg+52eq2gkaElzdnuzJyGeL8R4qlAJwNlyFiF0jph1TSdHJMTs1q5CbR7WF
3eupQWitLcSdpcJmy1A8UGPAAtCK3gOm9YclfZEW+LQKYYfSmspOmXALdlvCjkB9
7b6QbZMefzChW7EeYsfcjvmnGZ7GVRZu2r9oMQZTgfd49cEMDxHqiZv37NpJLvPa
b9NIT5MXVXRheLnbxRO/Cyya4rm4sCFMo0pxyIYRPwSH7M8SWkv1OteC4i6ylCyg
rZgzzr21bG+JVON8cfjWPD4dAfLKc74bCp1K04GL9ARurN47TnnGmESyPMeOv0Io
redKiYov67FQ1QEUnX8ApeADkBdMAWdbuVroUi59Sqzk/XXLqmn6LrQeHdbTeal8
lmuyIW9clQnb3W66M6i69GbPXXYPiwpUHxPsylJ3l7DChON1wojdQPrPIoiwUbFg
bM7vDpiur3R9vQ474EprM7VcBnrQSaVfQ4kV0LhwUCLKzYphRsc/7DuxsxSAgS3D
TGDj4WWjhSz5Eu89qdgj3gL50BYbwCGSWd7muPpCZitZCa3AqdEhDHhnerOjBtq3
Rfd/uqH2Gayvy9euKj2bcFVe3lkiKNgt/8cwi6TQ5BE8mzVDvcR3VMaI3yWzBWUr
ZXAQOYIaZ5FNWPIOH3KiJB5pPpjJisL/BLC28qgKuUnv/wD2qRjQaxCByUnlNigA
JoAGny+0+jpTGsCdG+krc1ZRbCxcyudLK8RfUGfTR/X8ME9PD8QKTM/KuEtvrg+h
IAfBNS4saj1JeUFjiHsn7VDVDsQ7sgH36Qo1RJuiWTamyO7N2GN2fPbgE0lZ5Hvc
hpSTejE9d7xC/wrxH+LbBE6Vr0rKgAtA94eHaFxaY2fUKrc9EP8BnGKBeccNUdba
6BAtoeAXV2b8jzR4W8RguokyBSZPMxQ7I1F4Wcgd9bSvgVyoT517yawS/BzGRat1
ISDffRq1LgVS1XXBw+TDXrZw6/SXnoGD7U0w9wO3yPxinm/p6R60oAteh1VXgUq7
hbvLWqEYRFuKJkZpLWLoYrIUH92uzDVgiYMD2UrBNtotKBfR+ToQdnXIfCGJlYO3
/WaREYE628iVNYD88TmncE36wfxWNJU0sr7aWS6GpFLP5spjSS9slXHV0WOyynMp
qY/1ryxDnU0/SX0P+mwkjVFt7p73l5Qqkm2OTIBQf6QDWEx2yrfqgI35f/8y+Twu
XQgj42DJZDbYKOB3iWl6gsv/BUAaObMB+RcSGxVkskdcTN3eJUfGkSH6blpaOIwl
pX9PTaTxgNqVWwHxmtUGLTCldvNn9yLPMK6sksaAxeemVMbKtXNxJpL9a3t8R4vo
1kLLAYrYHHvKurGDshfF1u3RC0FP4jnnfAiiYlohDomfYnF3YwqLqf8zzOXp4/sX
909pv2Z2CfMDJ3/n3vgqvNvqV/rl+/177X+s7uBIaxNUmBqZ3rm6GyXKdh+E8lrK
14u1FLcEBqP4KWQujJPa2XEDRFs1vR2nSMEw9XABTgOHIiBGaL71Xb2GzqUcjV0q
kbQDNQRl/uf8UQJGJJV02ZSnxXbDv04LzNoTk8oTpegasFeyQ2nTT1Gzjt4bgE52
M1AkjlIQq8eGzn4/bI9zCFBXGJ9tcltb1o5QIuclBOUBPrOkHeW7b0x7WrezjuWP
NviM/D5n0lQDrIg050z+CINSkEslrL7/o/NeIJRG3LTsIWFSAKBvi5qi23gwnS2A
kEH0PD4hfnvDCPkAOk9c1HYARPjoyB8W1A3OrsgCAY0v9zX4GfLhzxEx23TUoaCA
OsCOMGwczJIMJzuQbytUM4BDee6M9eiaG/yaOcIyaf5Y+uUIUNO4GlQXzo7TLiyG
7CcLgGelramnMDbXwwEbfgVxGe5Wt0TOIw7s7sA6S6YRWbgEwM/RKofQBNaj5LfR
SMsHAWzwrY4uhJj4jMsoFWnrqE7i1qf8I9Fzu8MJb0LMCDwjZ6zHHV0K4+h3D8yt
APUEAhGtKGqW8fbtGfcapj+/ELjZOkiLoZ1GbfoRTkRFw4gI2Wk+OOHtQ1/bXeVA
vc7Egdo0zcs2f3panhVh64lJfxHX3d3o5mbCuFaSnVkNECAU0bJTQFFU/H90CVaR
/vrUIurTStH/ZzWOVbhHJqFDT7ThYWcWhqt+VM5L+kguSXUeHcfZLzIOfmUPLccB
UUZOO7PHcroHkmHdYOInqzya+Brt0Dla8x//AE49OxPefLGJYuYi7qBqjo9eV8PY
BHjIJ7WehKxRFpzar4K/GrB1f8S8Iov+Izv3VNGl/zWNj2Ovhkb8pqaqFDYMjrSM
htgNXNwVmmt/D10opGF7BzoTGvBUWIRtFGCnkAVBBDnRXnUM85Wj+UZZZI6W+CXE
oHB6goFpT+beK3/fvLr2WH2jCz3Dki4XpAyCCIORKs3Nu9GbLO25g9GUjuoZMGAy
7RBp0PRkyqn8J3ZoMQQGTIIWXmRxisDBAphgUoYxoQecoCDELBsBejt1Z4LgUfBV
BNXZBhBRYAHcNjlCjGrI7Adz8D1ksy4meXVbooTs0johG5kLcgHLDTLIDnYkeq90
9VGCDloNwMS0wzJIWzxc0gS40f1BXhxx+K5BXyPi+PjBAMhOTIPhWEjAE6PavkyQ
vGh9drm+fjaHUD8I6yHaKerrzHVvliC7B0cHAeAtgxgBDoLo8kssiFS6I12MEOH4
JarqrTC1RBnTtDgr0OnGoH2qmsi6ZhWblteWl2kUgTJmmb8a+DiMiFlqcLCocpfv
h6FoFlcskCJXCP9iOPliejTpAwTY8Ehsgfewb/MDfRAKr/ZAHdKbgxv6KF0YSZEv
PrxM7mcb8hf2EqPRA047hfkiuWXSXjmBaoyGbNXU8Zap68rpwWs7kpOxSq0Zx3zM
1Wi6P70CsW5KdHU7dDoEL8Z/7SXzxAJnUBbSuSvPP3gQAp/C+LZYFh1itk7/4UEF
SPuWGuUuZEHenl766hJ3uve3azXodR4wvtruXcnqXZ5xKzWmYw/l2Bq4WcLNvhcJ
uYBeGsuf45iV+EmgoWnawTb5G3TrIcxuoqgPZF54bphf7jkBaoUIJiBrwkdf7Tzl
tmDB6ixRr2OeHqx/8+F3hU5VdWA5CKOk/5t+WqzL74R575PhUQY+c7AF25/yx/vT
NuM889BzOC0wN9kHO4FpehRFZ7QcLK+E0c9W9snk32lIfnwKafaTZs50DyOHte9N
bIHA3ww71uJwZWCgPHAOgTQIxDVBo2PNChlGNnz7EZzlzLAMNqh1yxelrnwCIALI
YUoigPMALVhnV6NkxYdVRRv1xSL7sMW0BSKUyRVCqAm+KGSnKa3m8BuHDBqsdirz
GfRH3DAcbK//On03qwCwwaXDdAgPiBjuw4y3D1pkXyosOMpr2la+w6dcwqYGYsIQ
6VPtqalB9CAq2XbTxfycNprlDBSWanvUrDUqzD80rhCRFEXvKK3FeGHebSzK4Z3j
P1u0CCIgEAtq3dRpGUpHJ0zAWReAnmWKeUMaH8bPKnebrw4l9PA2d8NCGZoF0BNp
60JdkVSX0mpW8Oa3OvXS8O0E21TL+yY14V5eSYFMUO6bqTDMb+2gAwpadEbrsFKa
pHg+ejqe2fzSRa9G/5KY1sjnUvJLgFLd7gro6kRJU9fIhuw/hCmzVfzjbQ5r86Bo
UtAx/IFuVA3gqJ9vvIgqC1LtbexeGQdATJa/fEO6uoBnL8iJSsKCAfbjMADJ089p
nMVoSZNWmAkfvGy9zFusxxjl85We4KiFU3gopV1Ns5tjsS87/Qhmkc+6Iq1Gcb+r
aNLHG77zP+vjrR0IfgSprPF8qLcBVUNd4Xv8v03t04cNQVCQFKWNt/EloDsjnw9U
wiHDtN/J/b7qBT2uSOcEJgsujDLdgZRcBr3juLUqgWxR3+q1eRmgoWgF9v9DFtPk
1XsMEigwqbDm2Ra+rzQM28bDe2eGwwaml2pl+A//pts8LQgwiW0XOHX3awnuWEOF
/pp/Uyqr0dhJ9zr/4VfX3bseAXixTuLKKxeB5GS2qDhyARlU64wiSnke9cl/YEMA
M9MxkeBjYGKoWBrS3tx6D/eJBOPnYylDRSJRBrIpush9eI61Jp+UY/cDgNCrbxsk
7l4EDXbGsuYtpkKwi7S3s9QyY+OuGet3Ie7u3HUrm5stpAnVt1TZYM3epS23fOV5
KrKrvu+Jnb9QRZ1NEeclRg8Czzep4OkQwb/mhHrCgXw3V1y2n5P5/8cPWICKLom7
PX63Lje7uOMMSkevQe0+q4mIs0MtOIDBH+qY8fiDzu5jnxFRLdF4hmUJQbS6RKc+
NPkSW7zRFIre90/2eB6h5Y+H/xyGfK4yyL/ebWByjUorB1aUZdLHrbc79roaUkv+
yq6xa9tix7VM/1cL8aKQKpMTPR2l5nK2fdT2ZVyqrrhKh863JE7SvOsQEIp/TatY
7b0dV5sVmJx6M5FtMLFHrL9UobewQsPw2d7hARW4v+O/64niWWiwFEFqXCcssaNR
f4mZ8Hx21G82xconXtoyFoLXJ9MLAUgyvqFyTjeNa5qnSMg/fMLZP49edkU8KDqA
oKwyFN60QBzRb6n0Wl4GbK0AqY0hQqxon5R6tZ1pWhxnBoUsTyWgFMdE0zCVrvZ6
smslitwOmGQyfcxuzY5Ht/MKqdf4Eo1th8Oy3uvWHB0J4PWRWrGBIzas/XCDE6QW
VNT2kMcY+tBpwwwJDNNGazitoOqhkGiPnjl41809QCU+qMRvVk5JESS2Fla4kZsu
6UuLWz34mHd/AY3DKw+gRAqBkXXuLaU7pUE4SDt1zjeqa9xQ3NxAth1BH4ef8TKo
IzMw6JaqLBl0wEk6WQclz1SkZGe0U1c7GiQTHB+XiqI6C1zu3B1ATOMahuEwbPoW
hgOIAAxGE8VKorUUr5AzFu97dTyrJhfnYekAWJvLhGlnkWrs5EgaxJmtmFRGVEV0
CMZsS/e7ViaaZ/fttgtIf8W5tlqBG34mXBJsZgFs7iz2d7imi97tH/ePwL6cGG4y
39Eh2qk35ZTkog7FBegXPs6hYezfDRkFqmX+tXrg3MVlEXuizG5R48xhhXaU/d5h
tkluD+OvXlzATitE9e6s1mhUO27+B5CHxIuozANnKz2Y7fnlG6BH8T7gbkWToXlZ
tJay1vleRYuG4daJtTXxOHFnvrwG+HZN6NGvwy11ah25oMjWT7OQljonG8qVNwjs
3837M/iRvrW7/a247sr+CQOP/aR6mt3SPeyh9iYgF8S3fSkO0if5eUcqD8Gh25fz
65i584K4NOwxrSl5dql1hfw0VseMyAj77r9YabdqWoWDDwpXHlqgt51e3UW1NEY+
LzSu8PrHgRv6Gr85wRCun/WroeqUNQQT082aIO7Mysk08H2h9nYWCPWSOZuYx8+/
iuopPXi4sQjYNI7Y9g1vJWjCCrgFrd2kGfcPHRBUReyC+nOI7j+TazTPYgizLAGl
fISpSTjNge5zSg7YlkQCJ0xusS9FOjqB2l9JXcKINqIJ0lZK882GYZAyT6+S5vTG
ncIAgVVP/5BtVRjfxgNYLM7ZreftGFzBL2nYMGZgOMMAcSFfOS1nk345/GFKxdVk
y+LJdusw5LTDFiblgDGu5z/iF7FPKDXoA1DjA7Hs3tIivbqwbgtyd3WDVyFDo0WQ
TOfMf7d1hi7luYRTLr71uLIYicK8kS0m97tY9+PB8SgtGe0ryzn9Dd/h/T2fnkfQ
lpihFi5RUPsLwuyoZ2GZgAY9q+0skJ7Mwq7UqVfOCSKFtkx45xBgDmWYKY0abB3U
qQ7nVAOcxQQCFuuZW/Ncz65tlpky3rXP500y23mCKo9uefCWK+PIrl9+C2l35FAT
VQP2V61qrffVxbwCFJFbZGWSDVCn19tjZQacMzki7+pUNQ0e+ByrQC4F/oy/B9bm
VHyoTIzKH+uZuXyUdBlWXJe1PVklCc+2SyWoToET6v+Hw/BRwYiLXJSrSMswfPR+
dqgQY45AdN2qTkwxLlR3zjf/DqaKModoiheY/Vtn5pxGMZUEb/Zd6OE2xbCkkjZk
YVlDdfov7oRNryyVIGL7trQCP6gHsbhre2rckdpAIdo+uMPbbzF/8DZIiPNBHxaY
sBX8jW9n2iCaQqmB2z0o/wFk9qtftHIexzEmj3mDcPDxXJHWhYH9pj1Mh56vRT3g
BHHbwo+2T/IgAEvJx8jqJG96kAQvdcRn770jeF7Iu2AafdCbj2dYVRt8oZpu97BI
XYj05TmUFg7SL24V2mIkrgyJIdnUf/R2GGx6zq6fQBB4OUFrkQsZ6HUXo63o3DaL
IHUSlzFTBqDk5jwm439yHakGgoO/NSAJ4v7v9jEhKFDzZvaB085+liqbdNI6jedb
h2SdS7bGYAcaVNFYJthdw+AE78tZZrqKfsPVcsakYIA/KdzuLjSeDAYemSWPuYB6
Jez6hO7zkU+eM73h/rBppwAvYJvMu4kyUEN5zIQJidV7ex/7ZSwncKe+hNmGVvNW
kFS9OsbnjM5b/Wz5a2YvsJ7cki2dnv0zxtXt/LoJFkeroGWZ/U/5r7BISmaUmyY4
lhgPo+xdnPz7yqTTch2wPQAJlsQE6WgZr+UAQXb6PwizyaJzQgXaoonFxRFXRkT4
Uhvf9zCIkJNXN+1Dh++gjAv485Vfxl3hBRSpzTlsk3YrjoxRrLHZQ1vw7I/h/Zl/
9qiHU8jfNd6upJpuVOWDCK0hduCIv/+kXn5+ZDBqKUCIPNIbNfK861XuPVl0XlY4
LMa1wwxQ7tlz1rlJucwM64PFb6Y2FQMtgr2vGFcGeQ1OQybyoVEEfMFxqNfSet7a
7dcN5U52rRo90C2Q1rovSrsHoEO+0f+j8gtaBX3RcJ4Cptm4Z/AzegxqUzP+Cm2y
8kQhwY0+cj7rmDSQ5/MinvvhEGbjPER3z7ton+qlKWm2WIrYpvWmoUJvnvkYd2Pk
p2QlLAwhBWqClDOb7rBYWlxeJTWgo1nL/bYtJKpVZdcRTPqK9+vfhXaZH+bFwBvM
9TGrF+RwVNOHrg66zP1WaeatAJkMvubbg3VUfMYAwnBgHoZ3sFvrycyqG+thq1rg
bFC5CqWWSNN4PHvHCHlrjuvFVoKILb870hTIDBtp2Wchb+SybCPBFFbVqGLQV4xa
hIyhCKrQ8XjahX0tVdPRKKVhvoYAoyUzT3a1ISvV/C0cyAkEPbukpsHDASOWhdHh
LJJTQaYqIgSyZtXhCoMSLGKWEGZlUEQK+RYHC7RDFnNemfz2QwD210FUX6NiYhbJ
ByUUKs9rugEc+esZNH975jXorqMHmdgnrbsn7uFDfLAYKyDWajMMQi6Ah0u8JYym
E4/M4Xai7wo9/O1iNkN3aqYk6/TDILr6+auG1gWSn+NRdVzWRSY2k2pwH2epX7vv
m3Remjx3hV0VR1tpzUMu1517342PXtqd/Q/ABQcmkk0olOVv/Zn+m+KR2Itozk0E
cizsBSDIPO8s+maKUrHecWrduOrz37i3p6Obh4co2OSSKTk0SMbMPfwqmtHxWj57
aej9pY8IyGP7A4MPopz5zGBpcPjziP5lgeydkvtjHNQMPtH2iirsFBWkG80xe9SV
tzSyqK6JN8AHOM1VtkklD+6q955RxcFWTE2XT1KnhRVmO9toucmgHJ5CBLXHexyP
G2pa06YM3j5GA9cNT71K185hexr67T4Nr0OcNPPmnuTp6YhSeWIMB5phJ+8eVPYK
nXTYoLat542+NuIRvUvOYw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
U2xCuzK1vQ6Deud3S+cTAoWnEzrHz4g83E9HCQBBJrQtsUFyKEOuz8xk1SUAA0sr
CT4BgJvtI7VeWYUZj4KAHH9hnmOtJnaCt/XYGqD+WKWKyavdrnLm4MI2EjnP8lZo
uRy5vniTi+Cg1iJof+muFOAur+gp3FCvC5xoHJWKL5npIuMhbm71qEvjTJv58wCc
wuPpEO9NFlnnm3tGZ2KjLFQ6R0tUWGpTk+9hINcnJ4VGjiBh6mxZhRKakozwJe3s
O7sXT3cRIIbTbvdlpVO7xz+O2ckcGXRP05mpGUXeUe0ViaDhww/3QN5oU0dfHjlc
NZmPNACV3ahXPvHP1Hrkrw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6336 )
`pragma protect data_block
trowaXkVwZcdHngF2z31eut7YPvMi8ejXfUCpSLP7bCEx3l0CGDxhaFQSLRpraNy
21r1buKRkhU/0aD0azLr0yg/cdivmvCoBh7a4iwkJTMAPuwBXOqwagEOBY0a/ohV
hTYsWHGphLUaCwUDeDoWMUmUknlnzQgqRgQrlEOymCHx5Ou32PdvyMEGz5n8A6IA
CX5lSeuH1TOn5Mmt0DtLdb2FRyJV9worXAXjWFP9zA2n1I4aMfSWH/iS0lXFPVCn
+Lw9CAP2pd+GlGnEmX0mESTNDF3XAhHRsZHrctGiuRzU1kbFTa7dohdzEPfECUlL
UqzjACRmy12itTKc9AkhWg1EeaAgMaBrMttf48DQltv+6yRcXx504EvZ/NB/K1ru
uASNn1UYNVu7Rils/BvQgTfUoz1ZtSBAOqe9aATPIrYz08/nmVnTSri97us707le
nS0o89XVKnGktv/rL5TUIeSfLPw9akTk/URgupkMYV7/eUaby53IzVW0O7FbQa1O
fn2t0MnEVmZ5GB7f4wMVQrWE5dvdcGVOiDd7m/mvUGb3LLnRmPwocWCNcT/HIPpI
rXrhcA48G4uzvuW89IS4yKszERJvOns1q8sjKHSuiEO5PZYCYD0yVNVN5gU3iIdj
GUbUBweUDvhDH/7t53gcRuQzwWom2RImN1taZYIKkS9xRB1i2V0TU3lqOGLLRIbq
wK+6eInrwOyuU8/6wH32hVN8LKEVSzmpNuQi3qefZG08EvCxLwy0npCaNnmxdBxq
ETHMYuo8eWTqxcdVGB83C/De2Mb9C3BoXNbZq+XCwG/n/mfjvTj763Ii6oRdqe6q
yT7LmuZxPk98DPIVZVVJ0gmV3iknbquSDbXsmX0xKNFBWThZj9uUW5cCrJOeHia0
eLNpmpdvTklJl6V5sI0XGmQjTf+AeCJc0FjQDceQVOZHl0LB2RhxL5TZ+qm7l/KQ
xst4yEtl+WZubPxw97igjqCxbhjibqqLuU3FAFdoakcnIo7h+ph34HQ9cci4lXCw
XKH4s3EBRmBIZMf3dytRaTRpMb50QwGewAkvSjpzwWSLvu7RUCkqctZbiLB8NTi9
DQBi4JpZHeeUGOKQOzUmzNAHedcZGPsaHWaG4/4gNB4lTmdaGv9LrT0pFzVrp/yp
bNg3aPAUxCjVeNYQlC2I4hTYqzMAEbZ4ZQzoqewgiUzfP2mTqNhIf6jo3dtWkOOW
x9Q5K1u7rEAAUqENv+qRNtrmssb1SPNI3sFAygmxwNZk6tRUdUoJupf85e0Gn38E
aoLGbv3SDZiMsLSdDLoD6WtlpSTTmJxOVb3pzYqm3TNG8+tAFrzpc2j5GgoBI3SN
/VW9Dq/csF4jtuVaE1Npiwr6HiH99L/qJmQ5K5FZboK9vAyVVOHs5Uq89ZhXNoHM
OFh4WrmVdTafAnfoeJwVIjx3JvALC/ulO7tXl9mX2ijOvqiBa0PbWkO5Ql4xSC06
tKwPJuNcT8gXwtErHQU6Z0RU1/3cwDvXi5WYt7Mtn4oiVl1ANaM71H5rpmsP7KI9
3XhMUG2CdsNTbiYYwd/hM4oW9C7kSJ0aIXKXVKWJAM3pGD0WYqBK+K0mgcalXHVC
YFf/2NK8/lw5ombB3vtedRAH1tTOgi7K+tELv0hyfpoi6kAdmyUz+a6apkGW88U6
34b2DO1jMhJyEGQACqVrVackCjyQlM0Bw4K9QagFtl0eRfxzqb4FVSFtRWv8EW96
hCb1CQouGtvYcgNAuqoUPf4g03cGtgp/1N2knf/Qf7xY4tS+rbrNxde5BzHlQdSW
V7rsU4q6iNvDKYfjNAA3jtSF5tDOy82vfjVzX16J0mjnGkyrRQPiow05US7vgwcH
Gh7Qvx1s1t30YMxNxXzxYh3bkOtvmsSLp39OSv4X+4zoc1vTNZajeojFzvaBBt4/
Wkr+x5o5egM8dTGovdDu0pf5qDMYmhvLXXbVcHPAtO5VrFhYHTNV52A7WOM30KTE
IAwZHMKGZXQBx8tUTUcnONAo2o+5sc/T/nXo5AizbKuJKJ1wUasBYg7N9VS1Ju09
20S9YFi2Br4mgadb6eEJJwHkpziAaZ6dMNnJxD9F8GWoB/uIR9weck5bdLayIPvH
QTTFiiAJKwi6zjGL1OxburdPI41wsPeKHsHp3S+XiMfB2V3D/tGmlZQjUzFqdUt8
VdMz0ECd+iiAOQfgAbALxspyLFwNk52vZJZ2k8n8hhPJbgCp3Ah0S5pb1p1kjhkq
SDsatkYjlYpxpVmMIhwA12wCIWQv7yLnAxAtZ3tL82/T2yCk4eng+v9jZGekiCam
+wFLQmYLsE3AeVqr7MzYnUeta99RjqYtuveMU2xLVBhycGrXGinnXck21BGyswc+
0HDl9d+syuzLPHqVZRVFspnOtBwYek3gJF/2GhL9h9wdl32A3I+NvYiF9ixHdtBa
24yWvz2A27jtCPaTlUW+19MlF+LtsqhLmsfj9SYMECD5bD0ycpDr2/PFTMdcFDal
xFQSiHllNZG7rK/I67qTgYEZMRn8sJZl5BQWb+PlyLrcWWxGgtb19fbxt3UWZ+mF
z5elpM8qygixYqNgWDa4HlfepEDONQDf6qvh0efpiLpW5Q3Wy6/2T6NFcITLtYT6
tqtMAC2CWUAhDQk5PBC3BDFcsCKChgkgIG1hW1u5x02rYr9k40ONt00rP1OHZssF
QfBxt2ajPWZI0A8GvsrmhD4mSjG18EpDxyLNrbko8p4Q3ICOyZ655bdv17rcnAae
jex3smci+alIyxjzdpvoSnzuevVxYHnXlmwjqVcou3yHqKP5EICaRTkOwvDT4V5T
tYlpyOqh34WUJaMu/T6mTWTBlwJJFEbCHhNaStrhYqoY+cV8SqS3WhJb81t2yrC2
mpJetFS7CC+R2qyf3d2dJoVasxZaUzzhsj/ybCroQdwDBSOUo192yR4VHgRvMb2r
WDnC0WNn8Jdlp0/o+HtAtG9pTT63fksl4XYTSPD9mC5+vij8Mn3ZsE0r4VuV2vVX
NkHHR0eTSKgbBjE5cEqyUeokS3MywyDrZvLGIcZs1MWkKhWZaumCmAPZO53xnd2D
KcznQqvmqXmvkP7RBNI15M8mBw7B7/LREgNFkpFzi5Tw6EnNIWjg2sm0lcjTQQUs
rVugj7vN/pemdjovGuY8Hm93dekIOK4ompUotpSR8YLTKgkci10gHLiWMgweNx8N
QZNncB2zuTNfJwOABbBO4DaYZLELpxeP8aDFyyoGyM8B/ghVB0RwrM5w9zxPmM9V
fTYnXIODHwUjFaLAWt/e1pL1pq0QmCp+Ni+cpkgenZ6gbFcTXmnTJQQSBEQaeojc
fiz3iIiu5Yk1JzXpruZFoYkPv8KPdNPdh5STknQE6Jm3dnLTwrGqzosZL0pVAWIf
rys1K2BF2XFHoZRDWjAB8aw8XLSHJlRu7W6lwl9STdaaY9syeg9GY+/dcuvca032
oX0L2Ysf/p7QuIzgFxpW8XNqLx7/V2siqvPXeo0vtZFwu4nTWUIXi90uWf9MYTbU
7/ZC6ekQ9peM9Ix3AFfW+VR/X5J8p8YtlEsYJLyyENoAJqbCEmbXWDNLmp3GMaIV
2h89jRmcq1/dfN2GGgSFNah4iu9aU3mtMUkxWUAx3bYkzK17eTYFAv0Yf47wU9dl
WOvSaWOsk+ZVd5g3ADm9rtWnxzf1ccHu75KdaADjF/L7BJZ77Xav+9yNrssJOKpl
k39KoRcizNkLYpaIEUokGPNcbLaOU32BpFXxI3yHRZjyCJfO/aUkTIycZXfxTDlm
aHIQ/EyXYf3jM78t5LuRcHrZApuwsnu5bFwiMgcdwlTbqu35XDSdbhK6YZhiyp6x
ySA5eo4lKt2TXKRrUT+7yoYQOmOSFPHKwm+zzaguXw4nXkNW4CZaA1AGFRsLWZdG
nGSkSbfmclwhQqSxY1taZk21ntp0tF3GH1FI321ejrBIC5A1Ketdu4OM83wGBAER
KpArNEQgFdIkbswM9d66jJDCtD2rEfbpomQdH+J65P6jF4gVbOmJReK9PKdq1xDQ
583idjHl3ryawGbBmiUGTOyEpy8rccJ7Lx2pkUQ4w0yxdLZrfsQ0iOuDzmAO7PAI
HhM6NVPIVjH4FQVERast9/tM2hDD376sDDXNpvpmkZH0h8+/4tQIrFBy6eOTTW4n
9Yeb3UFwI2j+NGkvClh/CI3pY31RZFAoWAUrNkLSiOWVQuhi4hMqgSTHtra6pHzB
fe6QHmU+jN5pTFtfy4v8OqphZ6TBZpFksQ69uWvaVDgk+pcgXuoHCZVrRPTT4N88
YotQQSk5suq4ag/nBBZGR78CTmR1XsRfBj3DXSM90ov8MUp1HLCTdXxcJG1dyjBz
Eqn9iCjZpV6IbYhdvg/b/gcFZiD2Hv4AsueF7nQQ12+4YrswnTjyOkBTet8FXXfX
gQZXcaGlmadOM4R7JwDPHYs5F5nbyrydzmG+ysMWUAZ9o0M+jFgIBVAWzetAaBSU
rAczu/hQ+2c0H3XyuoOCkOsi+B5mp6l+Pd6HrrTxViJ3Xs6yIO+TJhweoYNXNAs2
+cA8YFjnS8KzRSoHReGAlt5D9SZ0EkQC8p9CRCECR704eF79SSCoG6YDwirJ0VU8
6GL7npBrFI5wn2aShZIMGJCingF44lJGo16ZzDRAVisWFRfgAWMzxtAEcJzyGF3T
GO9XDFjTKg5OXBM+PvHXYDMVKDsT7HZ91/gWlVWGG8mYeiysQL949gfRb1rWq2Po
VikMahWlXPOeEWCtz8zAy72ygx9MisCbt+TJyayLe5JMqJ7QU+eHeHInkw76d3bD
49cTRmT6eGboLBr8jr8R4TTvxUYyZhCIyF3AbYjbzkePz3rejMHslIm7NRIPbaph
zX3of2flOXbYRaGqE1KjndDNEhjmIdM+zNpOE9KNDHexmPZ61fghsXyYB8hFBwtP
vsYiSYQqNKFgf4L89pFFpNsD8KrlWChecpBaUApIDPq1TgdJF0lxrcQItw6tKqpp
LINQaPseyqbtlUKGaGSswP2ZGBx+tng0FH96JAWiDik4D3DJAyaBYYmyCle9+0gX
tOjH5o3bD3QKLRnDpwMpoYZVRJ11UKHgy6zI3nqHkwotc0WAqdniGm43RpEFRHXA
Y7vlKnbAWylTzxGCWaVp/yTNQraQyACPDmFqCqnb6RSSruQPXWAFe0iaHnO5TduR
vEgT606hRcI7SWIcPkND1NCOyiiwTAh8xV65Ndm5wvNU6G5yAw15EgYRleLSOqbX
1RDtnyBM/pMPLLK/fciEMgmdWKHBT/RvWJJLZUtxzo/tjzWaMqSs0zk13x9snMaJ
N+Q/FyhZzxZnlLJ/wZBJ1vxCdBzDjwSTZxyojXbncVoNkvH0lvdRKn3mDygr1l/y
+3hxNFibqVGyWOOZy1p3BGeMISHui8q1Y980FGE4G8LMLCnirVE4WbLRMJfRy2aS
ejk2HV7RGvtj7uIwIJcqEq/IdlSS8+E2QvPV576MDGUcbDxDQkRqZojaEOqJi/o8
aIxCZAndV4APjvtbx4a8Fyu9UJcXFg1qWVWw0uzfUUuzLRi12yUmSq1tKanYqeAF
JR4ULQEBCsTbDR2vw27h8xCOHr//ChnrrvjMV+Mr1p2HWtUmey57htpEHBxCv4Ey
sD1C7cDKh3ewutJtSr2hN+IhxHJJyuxnW3ALJhJqtS3/Ngwbkc873vC7Wo6R3cUj
+Mi3Dujz4wL7yEhhBjHDx14Q9JyvW4Q2z8iKYd6u/mwR9L3+zJtg4MqQNHiCOp7Z
xAcPfSVvgaVETmA3YmrI2eSAykz/lA91h5ivioqbFwnKs8LDe81Yyol4tFgETTts
8u/mmaTrfcr5dVvZuKNMUV3XALO8K2noBVDQS+Gfs2FDQXuCeii1WOaMa1e12Y+r
MoW6YPjCVcUcHWA0LFKpm/RY1cRqzRh97AJq+8K+kS0dtKQTwWXbgR6BfgVluC1F
tsb1ZHvATsMnvrQ4I6DMLCi/yfhIs7IbxdErWgH4vKmLscHsNGHbAoruUDiFxjiC
eX+V7qb9wFHs/RwRh4dxx3OFk0Lc6JgKj6oWnir11ioyMZd9DEf1X/4ePZIFgHYd
HgVpBY7mWQC8+X/UA1IUHNSX+P1A/XZ6pt3uEo6y6/t5oO3FfgE7TyHDg7ZFSgBF
pK+qV8bmzDw732VLSz6NUb/eo1ZaqedcFqg4qPAC4xuKdVEwDqT3aPUIJk06DTEZ
E/xL68vMZAVC3wurVupZzJjpdd4GMGlz1QxkiQAM5OrcVDTebs2lAEtuM5sIblBN
/TexGETjtj4pYE2biJ0z0MsYVoQX3TLctBF5DhZ1m5wE8Xj881eQ3XuIO+exq0B7
oVVW5yKqKMbmXj9axwRwxcelbGbFYsuEMs8JOjy4aEzVtVLn7XHLlqWx4jpHfkRd
UU4bfCZqcmReIhJcvqjBv0HM8mPmrKKKiveMYdiyGbCViQqzj35YvZqU14vkaGxR
nA3HSbgtiCJBa1AbNFtSxaXhG7oPqQPF1qwY9CWEkxeyIh+ZVH319CwZ5ixJZFLB
KIB8GGhEblchvqIOZm6TfTn/bILHN9DW90ECRwPaLEVqqMUS3rYNMK8wUyPU2Xa2
ZFq/ZKYTZ2kkife4+f7wtQ16qSqW6FHkWPfTFd+WgBnDCIIHlNuBfcp2P/lnXJoM
kJH53htlqF0SbsPdIA/PPZjXxOlx6iyHmCkc8dvPR3YACxdUKMSIwx4QGAUkbbac
2XqfrDuYaeS7t4suFIJqNL+N/IwoSmsc59JZJ/zo3EOb3jEru1vXzbvkb7t/OM3n
/F/cD5tJ27dvFOcXVmpdhm1QTB5d7f5y3JK8UUy+t0984WxKf8K/+guErVCegOaB
wZjOLzLTG4XmCOhpwUkS/Wnsmtbay86ibvYn1MO0U45iQGlimvCy9VeqU0FQUjKv
eGW4dKwR7W8uvbgqrIFLMEeZzro+rNfJmrcxT4yQk4112sVKbg64bG8eBfnhA5rp
W2m/ZGUbk8vmMWZkvW/b4DTosDlu2Cs+Tz38jC2z/L7W38jggE2xI0kt2S/RaObx
L/2uI89xPqngtoD2XV34744WcDKOBT5yuNF4Luxc4fiL4892lr4828fgvkUB7M41
3ZATGPuJED4RiBEWyXKWCM+2T//sAtvAkZhOZIwH4vNP43sGh8JnsEKzQauCbNeA
y4lcdFGTs8XPegbEYGEWF+vQlvkfE1/a0TjPDaCtarMQXAxhg7iYmaIEtNw2vWbx
ScfXWK2T9V0JjIi1cHLg881PN8uMIk5bU2UqE0aF4NqBjBClHH9mppfK60wRLe3C
TjXPBFqLx5+zYo8vicvEa3f2VF5R/VIXmcc7VMUdeAiSPhkMuOGXOqtKve2p7Bi+
L9h7KC5xnywLBU3j+i7CVT6KrMVLD8MC9HAaFDKOk2BCofhl5mU3FZOoduTm6758
Nex7I+r+YbrxK5GWMJWHEfCiNCbYJdw4vAD4fGnQ+9+33ebxYHvxQC9FYkCUQj+2
VXvqJk9mPZzouOGed6zoIyX2c/IjLYhLEsWRo9c3FFgV3xOz7r3nwTXiyZQD/GK8
QeA0SRZXi2C3ux2tUJf9RfP1uls5hHQNj9mcsMQGJruUEdmR2tE64whmB0Rfc40/
QvZRiEKwvnDSfqdwu18RblXCQ27Wg6E1SpxS4dc3fXLkQUnxALhNWHYtu4zYql8f
MLzVwCsiUwSIjgRhbLUK7a2mY5rTriVdBZXinP2HVJmJsnFmyiyx56rBk0f9w1vO
4jxfzX1eiIipAiPZA8mc1VuQSKtiMSqH0nycANgmf8qtG6pslOsYZz3k2cvyFy4Y
ymwAHy/Vzg/sMllm1AhXncob7CkkF6GuNE8M1Slz9DgCRe65q6TMfkRikO5p53e4
qHdPEntm+ZdpGooWNHnp9+LUOYmpNsl81WoDX0Hq/eWoL83vQeHN1xJkBp687Nes
wi9e4fdndvYtzmN9HdeYhKakpsj20Fb4tC2H7hHP1UdwSN542bwPZhPVWPXW5XJk
BI9LUvTJ7XusTC+Z0INOdx5u7ol+O+s6EMHp+9iCwhyEe05rifJrLVGQZPL3W9mJ
ghaTMi93rElOnGdKq83Ftuo1DL1QWUPhdhkK0OpuwR7Rg6nnROb2R9uobobSAYAf
+ZqUanqFtLH2kh+NeHC7RLzuuINxXrELsk/vW4tu1ijd/SOHVDvpLv/BfOcRgHs8
hTq1GW1a38cDctO/iexXQ/jTu1ReqIafvS006iHbSIJ9s8cmeF4F2+LE7yU+5++j
JYy/ks+Tcoy74HH2doNQQV6OT6FsDb8eI6Tzje3hXetLNEZB30DDrjPlIrHjOAMz
ZZx2LyPfGLATc63bCMu+cj/+4N/rfYNrJxzI24cEc6IjpvdlKsYvPlFi2/xpVLa7
XeC2UtK5G8UgfjKtX0FEBZJyJiMx8U9aNzt0FD+yjooZY//kktq5tsqcbHcalL1K
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LPgYtFCGwryBztmPlHz4/JhDN/Z6bHGVtHtDEfmw0eEZFLls64OId7FiLQqh/PEM
UAFrcqcnmtoYb17psTwIF1agJ9BzBhoVgqtfQfVxLKQXRad5Xy14Z5YWvwHKe2tj
gh8YxAGGUKKu4etz5MJmFgorAwxnCYwka6M0S44VMgYP1dMnS5w9Nz/bCEnRYZvM
d70LNva45oQYYfGBaPtvsk2pB9fCrQecPQ/plX/WvuqdXgIu4zIpHUPYTN8Dof3M
+017FHI2fyrKCwWg8+mjk2UtbeXkTc8fQ/E533U5SxsFS6Nrr7z2yAajOd92sFpd
DTAW8UlRaVs0eEyfNDaFiw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 832 )
`pragma protect data_block
KBn3xsNin9ClI0TBAzFJqAMgj7d2Se5FXHjiKrDXZeHYJhd5oDnpeDWcXA2GQ8ip
Y2h9W1WR07SHpDtO9shPcUP6onCpGr74ESmcf5et7ojRc2Tpxs29VuWhcwbtv/Zj
l7t3wRuMj8KO9HXNBzfbUCnARLhXwla7qtiZxia0nAnokv/jvLvH52ZMFC9NKHzo
w6SApbn/WaNQPPZ1RMDF8V7cY7gBmJG/soVbltLFt7QyjYOGwqsvUk2bN6bjbSSz
aEr47jGt1F09JGEBjyAVjK5aZm2CEfuQfMvHbOIAwe90Bg5fne3c9Nc3PUZo16vc
H8eHwp/AGfu5fsZqu+jmKdviKZ9slax41n/Obf7EQVsaIBnJoDB5/4FX0eGVnGFs
bwSQGhePzTeam674urTm+ZXXDjDKrTbvuSx31N/bw7SFXRBYAw8TGR/5rTXblWcG
Ur326dUAHtqQC09NWKn9OqoBRGmPGkL8h0ydJ6GUqC/eagiPbsKpEuZIpwDhVsi7
HEbYijlNgngJ4N4RAtQtsibkrLNUfVf+aGs8Vl42bgVoJNyLzxr8LgldPj/dY7yS
FHbjGNMi9IxnMQiEaQqvgm756XxZYu6MrJzeqIy09/UHjbXeyi3K2Ain+sOHUkyb
IclHQKyP5JmaA0DBSicCecyI6DLbU3S6hmg5NkSwPAHw10qAQU5x710eN3JEwIpc
kAQPztlL8oyGPT9nx0EGZdWRWRPiln+Tg4LkoRKkoJexOR2gwO+z5aotwQkqz3SG
jpq1PH5Z5lDjS9UQ9JJef5l5ZR7ixGkr8Jmqljq39KHFbdHCc2o+nLrlO/eVtk/v
/u90l5jdMVgOQFHtDSG8Ei6bWyml0eW5qd3QkImoXYk4rV11IPp3pcHq5FqHZ/jj
f57gHuu60kkpLElW0S1rhKrfzhv8bfdCdNFc5WXsrqdixa2QKB00u2VBKKO2XWNs
L4hQWSP9am0SZmASoy7J4+3C6LtOQKFl6SGMrEs9TURbdPhhWdDuREIe4xBhcGam
AyBXv6WLzijsz5L/CiDqhQFaTfXAmqk1DHH35BEgwAUZJMf1u4WNS3zP/ZZE4Flk
oeZeZoIWs7/EjTgE7PxdbA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lnCjTihtvfxtpwyniFuO4upuTXpLpGDBDASHury2f7rUqDvAgl7B/RjSA2StirG3
i5jDHOoWLXejs3ZZ0AUEyQVAb99KGpvJe7jWMY2U+NhVBBrOwAQ12oIWXcoNJqre
3GUqahdwmwnUUkioT5sRnVrQFy5dATM1yHcdr+CgTjuhbVmAV0arOhB1gLgqoCB6
xaTwHXDND0Ke062MyhuaNO4D02+KXoYOz/ZymFTti5A1SFA6rOxrIXdFfsJYAOkT
qqpmQ23M8ZFX3Dg6iA5wBoeUm657Txu0dZV2S1iCl/Y2bi37ILv+0D6OxCvJP+yP
DCO6FpsiRk+HU/7xEASOZg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14000 )
`pragma protect data_block
/TZvo5vp6q2ZZoM9k1VSfKpLBWBqXEa3a6qtJlSAwAXFXK4q6hdO0dxms0YJZ3tZ
G4vSNa8AtvesvY/fhD9acmJ7oh2pUvpgoz6PpnDmFjFRBDoH/JID+9vTXiv7d43U
xSAHpWsObaaIAUO42zmG3PtMNyF2Mob14BKt0Aic4o6ULMjAvP0PqSlezTrFRdD4
0LEmWhBcSSFL/Zb/2Pt7XCyRK/rh97axfSZxjlnStC/MIpZvEtWtAEManSmP1P9L
2SryPDEKp86OQAuWXjuTq97PVpWMxbr8+xeDBi5ilfWVPeGYWLSxpY8aojS/Yg+w
Y3Aduf+keeBEB5+1nqDSdM1Gf7NqcvPQseOPkassiN7VXDFuShFA9pv853Q0KvnQ
PiXMqzGuPuYtbVD+fHFJAw3YL1EHr62Xf/qGvYAFfdMmJangtS7WdogEzKFVQjI9
hLMSdob4tmFq9rXx9Cx5UQebXRqO139F+UGDE9mf5K3L7igdU5MiRENIlU4ZOF9W
zkiH8Tsa/5RBdyJ7FIwreMAKzkde++VJZ0iS2MiY4zTtHSxdEwR89lHUTI2DjWox
1q/QV798xebWSAzLSHeE/gvF50LAXsOpRWbbXjUWKgNRMiFeevmVaOerzYm93wic
ty3PqamP/WHTRbWsuKS3EFwYNSZ6C9Q0BhNpkV4VPneM+3yd32oPPmy/yjXt5RNJ
/VE5TOccRdeZFHwucMukoTKIpNdpByssg1ntG/YCP3iZbnCBEDHVUOIT2jodP26U
cqC8xK2VRv0USRRWfQdK1bVIvrTf5aaZtoqxKlDgrEL+1JrKwJAcOpLTIpowBm6N
s6cm6ApcJtZhvE6znmqeFvgu04ImWhWHny2RzYD3t5z/srA1tvbM6njyDX4l92Tj
iRa0C0fu8JWQJJUl3xKZ0yRUEEbGI5WQTcAM/SRqFJR7hnoAcLkaobE31vxCMYt0
xT5BEi+/fopxDAodswW2s/azMiYdTQQfHsibXbhpKz9BA2mD71ZuoD43Xik2jw8z
uvmVanpD5HmNrvpBxqA8+ifRv3dYKNLnoHy4z5bqG0a0YQ65A+cJ1ZhNxNeLcxSy
3x7llOyW0r+TDm+CalE7nnrF5lKpRXImG53p+zEurmPJht9MU+5LXrNcvBWr+9sU
cs/ySe8VaUlJcAaT4/LscHXGumsGuCOCMZLponl2yg0e2VjlRdwv8om0MZJHWz26
qlRi82n0HY0311HrefrjfwIOSswqqNQOMSkKwHHIdMWBDr5n2/b9B6vulg9uZepm
W7VImNKYqKyGQENqxBtCeqrOBChONbERTS7SgFgQGAtquvdAzILvBMfRdYiNZg+i
dYsDdIs2B6c4Jvr70FaFryuErfsBGkWRNbb+ItQNlkOCIWSiSxZdJKGcK0ln9/uR
ngDMCUbI2RFaw7tuOimm5xQRgG8GGJA3lOaESn2bl+pLE8LxDjenPNi6sRawF+Sa
fRut0RDJxHUKMxLTfyGonYQgj87x/DmwdFeqvsPEDIW0pdOt4fgDjXB1r4EYdh4L
h+ivbVkN0TOYKarZOPs1I2JQ1zJ5tkhFNHTLN9yN2HpwU36b7oowUyuU2nRPuZBI
5Ehzvo+y2TgSuW0v1cfua9JSE8e8ctdo7G7mcW3q5DFRGrlmAGqkrfEj8lB+ehqA
BliBIC9OdbDizlDMZ+uUNyGmR56YL2wSnwtXyl0c2veF5H58816B21rhOuOZcsIO
NTfXLDD05HhHmjA4+ppvTF7loz8roBMHUE2Xgj5QbGxXPMB/D6w6yjHf0MEyqBJb
ydcrl5hytKOslC0UyKQrq5sJGiEF0iHm+2wM9gAxmdPV3Nn8CQVFQ8TAO5MXesrc
VrECCrjcMK7OeIXJC1c6zYdwutF1FJQtq2X8+wHP97ejBViuyPtoDxmiZ2dv6wOu
sdh+gdbU9F42xvHZUpnRTHwdgmnpSzwiuUPVM/t8Va8yx7bu6rWgi6dUP1ZzdpQG
4YcfEV74corQ8wofgfgGGkmy2Fmzo26enUNcRPi5YwclLpgqQgWCNPTORBjyUs4o
Y+9xS50OMVRnbGujpPxmFtUk02SW/kioqbFw3hlcabcbhFWZ3jr7EoZCU2muI/P+
/V4LHqmh5Fzh2MFxZG/aWXXn+VViljFKbPTUuIzXVI9E/JW2cjCxzYhwmb14ChPc
FcD8O6YsUCuDYHqM+dCTf4vP6esKbFz3aXXMdy89HcpCUaAocUXGRpCRVMozU2Fs
5selLSZayqj70jt57sovMQORIEpe05UD7wpNTxG6qymDUjKG4oEumqs6xGRRLbUV
KTrIxGbKf0uO4oY/cl2hJrHRq0K1ueegtUpwhaPOXOR/XFImD9A1U6mJA1c1Ku1l
JaOZDOK6CtMcNh1b5yHaw8hlv36ZeK3vzcb43u1b3KGzTyTSuwwHPtSzO4trM3yu
lgVqj1oeRddm4Jc+iGa62wd/cbTidu/bcnoAaWskbNM9k9JzvHVaWPfIvmAC63nx
7qIwQmUYO29w6BKoCjPaqdFulaR8d8EHrFHDjHqY68wXDnSmPnJkUpc+8udFSpEv
OQIhMLHDR7SBnBlisTV0Ih2+zBNhGyxRMjCPuYMpm8Wo7d6Ouwp0zb3sPVtFJ6oK
tY6j2LZoK1cktn4oM8MrIttFFXt+vbtGTR1NybCqWQ0bHjgaTr1Mf3ttqiiuviq3
cggX6UpPWioTxWyld4qIumQwKn7vgruW7z2qq9aKMces6oUCYu8c5oYiHbjkrtMd
QGiwF3fxdOEmOJptWqhx+Ixsk2uftIv1hBQ4b4ZMOAytsy3FZLS+1t9MV1MXRTaI
Y/Ur9wLHuayF7YLfQju3Cdwma7NU6pAkqwQFkS9g4tz4mJRxNjEzxFEHFmq0IoUt
cMppAOsH95r7Zf9lqOVV5G0v7vR0MEj1dAOk03HFSR3u8ItpSjpsFdSd1ZDjbPlY
Pfbs6TMQdq3p1Gb8+6jVMmCuQeCm7YNFjfRMr7N5jm5sR3nO6eUgEk9MAQl4j4hU
jd2ZJyuaouC0VxU5TOp6H64nld/6WA5ZZENjIxzXpmmNSxSFQ35KYD6ZOOrIT6EY
Vex9HvdaP4LcbNNkt4ZYyPF4LIUoWTXN2qxfoEs+dPUmrz/be/uotpOfr9O7lmAv
mSKiAgxv9JXNIFPIYm9Fc8gCHQm7Q/XvJ87YTiFFk2e9Xb/JY9d7v+/oBgUVyfyF
2NZ7SgBgDmYoV8Glv/CxL3V8Q+Qrwo5ZNgFmGbNmQnR9+GWMEbMtn/EDjcroMLuk
FLfubd22++5xwSkS958fi0OLAMsASF+j5Arpm/tcsO9D5khpNlnziTCVEUffBKDw
7a49/QkhKDOWL2jz7hjvCM1lwUzsD3evazgA7UJCv+Fw7967sBIkaCfQapSgD5Cw
HnU3+nkPWaHShz3iIKf+qAOWzpm+xCEZBHcAq8gD9YNGM8k4cZbgHL6TnoqPjmTB
JgNZvaddt6eaSHqHRnjE6mmgrgG8FB3v6AeoomuizbykESpGL3Nxu60KO3s3Xqkc
JOFNONVS61YRieamAiGfY7+VFczBmAqrPVgKYVSRDQz0N4bkppkSHZgtIaH9IRUJ
60iFp9tdLIjx3kvOzBJUf7OXI0fqpt6+A7DOpibS52yeTNkFZ+yl2PEAtsr+F5et
QT4EpmJavwEJ6G75v4kyVgncY2hTBPcRiGG8F8htofJGPa35OwchnczaqQYNbiHQ
ZFKGGJGNLVRVKJEDrD1qlecH2R518/whiui8wQFjs4ELihGvS8HY78ExHhx58Zjx
ditek9wDR7AXepLGrNeqtAG2DAKbKqWZwl06a+W6PKoUjAQSYWixMl+nlVQFWFe8
ZL44qCqY7iEMN5pb0uIgCVzw3GeAmcNMKVh4f9ya+HShK4j6kkr8KHVyA3EuCbOO
AfvdngKSbIHIwNnCc0aiuphMpZtOQCNtZ8mtG318/5P0t26XSv6ynChw7FFbDAkM
NZsMI3ADdu5SL5AtcCP+nXq0+3JoYga5TBWOlo15649L5D7hMKE6sFkjs/mypZf9
JonPXObASJiANf+R/RHM5IC2A9hBsEN/nSAogGkJm8ImXMcjH4uLLqvcEX5saljw
q0m3qqrpp5gZyFlkXL2yUXIaU974NbpXIrR9SGQqo7/K+2CzfEHOw5GJfRhnZ1EK
BMcifbsea1H3BmRtwwS1c/Derm2V4BrFZQHSGG0C9mpcXJ4zAQ8zawRK23NMjRs4
OEPrs8miuTUSZow2GFzIsRk17xkUXAHTp2gcxFdh4h1RGXoH/W2GxWlKblvqDYJu
DdY/uRU2cHiLP8WH9gyCfRilzzVsIjNU3rhqLQ8vcXEYrat5jf/Gkyz9JfxoZtrc
Po+egU8it2VLENWlkIn8bIqQ5H947X8YWd8BqIEmuGWetril4Wp/QBiLmElIszTW
ZfQaim1Inqu/TFAvbuQiqCe/lam5le9xAl7dlXzysmeHi5vWyxKxkyuf3n2NSdmp
T3kJgoszkHzeVIM1hONzPHm5iZqYFJSYno9MEDaJpcxcYfX4jCCI8ZeflgsR2PDy
7kavulIjQ0zFyiTp+9qmlTzHIAcggJ/PzkY8CboR8lTDqAMAXyBozX4YenUXDrvb
wj6k7haTH9aNv7J8wsQREnkmTqYFwkuqKRtr9gswX2R1gU6aO2d727S+INnAaEBO
rzL6nqyWPAKvbdf1bpWyBMKS6kwJZHRwQ672fmSt4laPg2IvYl05tbI8rkfwoPd2
uL6sc0SnDY7Vn1BM8axNrYtt9AKB8tRSdsR/0t46T8uVNC7ejgEXsB7dBMzxmATe
9iMQjD0KFbePDR+uWGgnER49SEd12+MRS2+Qk6GzXRlM0YLFP7RKauo/Z3//GoAv
9ZPzarVIe/Nl/BxERdTTJ0v9FOL/W/97UyGZbWgi+bytaAVAGMYhXLEGnLPhIv3/
0ia3fzJBWk3zGPRXNlKNJM/m/0S/Cw8G458yrQSGd66PbMtG5/LFERDnkvwX0oND
dS5CJAjKCksG9xCYpFySoB11JgOE0XASBk/2ol6mbJMdXIJtYryaXAU33K7qgEZc
cXelSMPU98wl1m+df06E3eedcEvxnzrek/af3cAIzWfUORiNDOjIj6b8xQyzA9LZ
h83M77unmMCq620sHeKASiRmIl86A7NYdBG3Uhqzc12EkvRnsKQ/JkdOss3fqSNt
3YQ9ndOgL0CYwh+zB93MHlwFz+OZyPQnK9eD9jFjMu9PU4P8k4mihVSLiDM3sCG5
oHxqpwHfwTbOLm2uGL29MD8uX/QwtQnKJ4I0pJwYnrgmedMpQj0gF6KSDDxbgO+/
m++5WqPUdCmuHyDBMjQglogBY8incK1FVn7tFa/07ArS8apOukzNIK637oHzMesP
IX7FyvygUCPGCR4Va/n5q8I9NdEsVyPjjas0+2/zwC3reRJCI/1DQUv/FPRm1vLZ
eg4uJI+Sxzri+fGRgC5mBNwN/2UGyD1rY6smyPOHQADuM16yj+oUYhdMAXCwXPve
106AgVohV69fX/HZFjnp6Y5KNemXjjCIuCTdwm/fbW2+5YjUJ35PbEOX0DaxKp97
TPhXsK3x6o7QLKTS9Wabo92dnro3YdXcBYNvNC9szf3Q0XqLXNiU6KbEA3VXUsYT
lvU57JYnqjJJ36mg20Dh/hMgwg9TfRv5ieYMtktM2ELyVJzflFjHo8YKA8cz8Y+Q
tbz3lL6/wASxBkrBVRWKGVzL7ZSfT1b7SX2VkjDPOgxc0vSTlbWHu9dlIF9hpNow
zMN2LWxfnHZ9+/r0CYfn/gp3lC/iCU+aZU+XxnlvHgIXVMt74OgqfpHB1lX6HJ3O
/htKoqQH5rBvIA0kY2aiKO2gpvv6eMbxFafBHi4MILklHixEp+lAlgH6JBSuoJF9
WEzV2uN3huEIPLt3FcvToUEvlrvfvfjvj3kI5ALY0nyUCarz+HyRAF6i3NJmw+Pd
VeKF3xBhCDdoyL15OwxedpFDeHbNC+ZFwGQP0Du9FPq1OkVVYu1qE00KZ7oiz4r1
PWXzI/rNSa0X04bdra956/73w3Sx4gVAEdoxT7eLU+fGFh4vRPnB0oZoh6jX+c9P
/872oQhilTe25LUCEGdeBQqoBnKV1MufGGovSemPXXPjyNPnZOOtof45WH0aSlFY
Gh5rBYWwvCXKSmGKKAQLxjJeacW8UvArZqd//pDsi9aaBJ5AZ6wWGFLBbh+T3Fdw
MWo+95bzRYXcS+DZVV5+pO/D4G4i8zkZ27GFddkSavU+BjzDtDSBKE34T4bHxtoA
xX1NCwjiylF+LnmJeJHjZ7LzFKEPD6ugwaXzAtJ4eLPXMzxVT0U4a1UVV5cDaQ8f
Oe4h3siytytt0VxFs9QfCm7rSoVVJZq6d8PCPFlD9sq73tRgM9AVY2FmX9O4X0zT
FP3zJyt8QYGbFmZbWsmBfleW7Hw1MqX2tzBtVAz5hYvhXsiNoPjOk5GioHBsHjiH
vqcPhzzSuvOqI9z+YNbb4MnqCYleKu79+pJX7UGWjkn0Yc6b2018xj8WcBSrg8Vf
IFlSM5Nb3LroHrhgRFD3e60fWBAPGwUVvsOCNOQBbdrLimCFT8U7kP8OoRPkHaiK
XamuG792HKR7ZZzOumc95v6wC+Up1XxtmNuW3T22g/StKhyQs8hRvKJYsgahSEvl
M/XyWzM2QCFUyQzV/pQ3N2Oz3DeNs/TtJJbOJYjL+lNZnLnxH5AbrG9ELvPdnCRS
x6Fd0mVXTc4f+NMMBA5SWI3x4jo3oJLRjf515OtU6vxZQfiVai+EAdqXEianA4UR
V7Y7tpgYF8VZoWxdAeCcqkdHbkER/1KddJTIckOnCWG8HUQpJ9TsBupzFczFXfY+
QOcgHOXs1uMXSur6YQgUyuD3/7OhwCBbRQvLUidMYCdLar2tZ6A6zQW4FXGWuKeA
Y1lz+TSbyTmWAvECwQwMiFlq8WBYreTHiGl/fAvJACv2O4qpdgOrY/kyRiJwVWGM
0juXSMJftPX33U8ZnOEQ0dVASJdFF1/o5jGpO4b4VGf5JJUIa8vFFmlXmpFOb2iC
rK13c99oQaXZEJNFr3PLZD8+kNr0oHyx6Dc3PUmlylNW60Eox1o7c1MwhKTTdKNL
M4/F0QqMuoiErR+bpEiof/I4QEKGPoELQtPUaOdnUZv7mZSA6/fTnoVhnfzxYvkc
3mMWO6sjEtkOl7JuOyrnho6AksK1K9OFPTMzReOa7GnaC8YS5r5/4WmtMG8KqIw0
XDJIrjnPOQvaKQCkUiykF0pFlaONF1/lJpgwU0Qe0S52UNEiwzoaIIk+vDfAPU79
FL/9F3+kLa1lqXyhmOCT3D1SvLPg4sjr1UVmsL8kJqhntkBwG8QXH/42d8CPQRB/
7M/dBfagTexXYYz0oyPo8or63Pc1skdenm06148wyyBUteu7fzgQF+YY53M6pWY/
W23VkBtkIBQzLrMNs+UCz0qSIlIRtqr8pA8U5L/XHXL1X9jKnoSTuE1xuqks37M2
dDew8czkGwcpDZOLxyFLVuER6+YkIH120gHSVizZfk/aQy4ervj7AL5A/NRPT9Wb
o8CQmVo13yHcuvi20Tn31T6HL0HX5wvNwK8LL1RBOMBF3tE4l6DBzkZHvYv5uYx4
uoZpELEJ/SkbplNZ1QjauK6QlDEPx+rpJ4FlJSATUxwp8ztwoMwcGIE7L64qxdVL
i54JPRw3hJDpcdeHUrk0SGHTKZb5HdSnrNCyWY4XX+pqaijPevP8NTl+lYMny/2g
3420dbLqNyBL+uKjDMUGJi7LxQbB36wRHGGT8zK+46zeUA1XpQ0lIvGwIJW2RM0K
I11eqabgb0H09GB2hL/MGUgYwif6uYtlfXlitbPPfEVxNpLCdqVJ3Pp7Z10ohI+H
HA6yxSpBLaXO5uS4Y47mp5UCsQTwy9DCN8R2MppF9Yw0g22RCQsc2KQ4jq6TLGBU
8Vqg5suNdomR7dPLhJgYDJYY3WcgU7s5a2dvo+CKfLCgThmueOr2pWEDbOGMX3TH
5m30pSa7uDYFLQB+nb6UCGA8ZSie4TfS+SrMyKxLh1vAgDbX3eYOl0GUdEiSy09I
wHBqnfNqC+UEzRIm2bkdA3tdkRe40gGpoLgddJ6/+qPm/xyk0yhLkP2b+KQ+KZat
AeBgp0tOcYesVr23i/kA2buOaxLMK1NJ+F+yGa12Pr7qxRtg1P0h3dtOvp2GnJjb
nWaMHolbhV/KgMxi30u1zklh3jXRJ3sAWM5SPgyuknS+7cgKfxQaYHbXrrWIqyaG
HS5kIKwh6Iz0M31hnNiroLy1QolAT61QUsJxaVNkHoO0SiGMxiG2HtacNOUWjlfi
JYfxm7Wy0h1PNpLKdsG8tSZm5//4OalNhVpVZH4ujcHSYarinfTqmfVAXjm88ek2
lHm6YRPH9CABYSF2HG9tiF83f8MwOvrNzIwdlwELzfZR5eZ/5ayfyJ6nTNtGbhjo
7uLV7woD2kQ6QmiJVJfcrr2BfEDJ5UP8C8SJQ/BfC1cFE90YMXIFD3P/AvkruifY
C+kKZHuj4aXQE5upAuQtKEo+h1UZGVQFeTegJk1jqjfbn3TEepheq0jYp+oyHgzs
JDLzc4Em+IQId8LHb4ktRrYGMHKkSwHcd7hoTsSWg9QTs7CrbmCe2QorcvE+pYNK
bf8xrvGruXUv7YWY+hHIra4htNDVVMHQ0HNf3EYon+0SVZ1Sbm2Av1IwOengPBA8
XeWszRImHRWjviXGQbntJZZKVOCQHO2j7sdl8/o+se7qh96x01QN2K1T/4paIzvb
EaFjXmZgE2B+MT7yMC/bumGOn9L9aaaYYJq4B5JyrzKgfrYlb2k3q3pMzG8rQTz5
k3GUltWrMfhfbAUcTX93ymMRhIUD//Kq7V3n0zczYs85Xu2NvjyDheabtgMoTks7
kXiC9pvwGCR7xD+dqRnCm16EGitNPXTl2yaEAihZr/wf2omhnOQPltFYE+510uQL
zkR0jpxn5O+IdVVCzesacJFyKWR4axAW/jTdhWrvm77Ic1ouoAw4j/YOWE/AQxuc
fzO+zg7/8q7upp+hXGSSXPtPV3Q5MkVVunCH1r/DY+uh/+oi0UgzfHgBQZOIpiJN
KElEYW8JJDL9/+ZGYETSgF1Vmgx+yFqpWnhmyh7f+TZnjpHZynFdqtWddSzNA573
IRGQ9gKwOaBnUfgXbdPxiD1TfdY2BZsMUOAFMvUrzwGJKtCf3fw6R2PdOgVfy1TV
xSWxf81K3q024TMOIwy7gnDEhecGtIzgcU6LgaJ07OTEuokTFvqmgb55zaXf9HIM
A4qnbAAWkgJusGHnuos0CRBVY2uYeNxT2/LRl7AmYDC6xRV9gHZKj21HpgZEEDNf
pJwHZ0IZt7BvxCkJwjOLFypnDOE8Q4tShL5NtVK1Z/1ZPcZry5rh65fE6seBLMSH
F84+qqkGG/CxYLvboDRoPe3YP6DK3jXZzmplqgO+khrkdv50nlLJ3ZwZKCYUJzfl
1hRtLdXoxTrzybXdELOIgMV6BrKIWGVrlTWt+UOqyI8H/Q65CapPMtV20v3L4sJt
X/XhiY45rXq/8EJIrpICkhW4MPxPwI5RI1GAnpkpmyQ1YS/kgGLLoAeg4mJtWxeG
vPw9TWuCFfx5yZpIRlwjMAp5aYiiEzzflPrKKao3dYIMqkxLKoobiI4Pc9HR+BWp
+VhKuWTFSUs7jQnl/HRkiLYE+hSNRBt8Z0CbniE7o/BWL467T+KAwOvyzusrM+WR
jKQWbvLnfi/t8xrROIGUWj9SXBOHtRUZXebSMMFapPEFolNOm1P/YKtTsBU7ch5v
pIaMXboSgWjHs9qfcPA+3Jvedx8C/wtQjXnE6Gw8JiTvhcjT6XFLubf+/FgTe6wI
QOi5PzxL2w43hGVMqgZtUZnzo98B4FJ5UPqv2iCczzcutBNErUPw6XEtf+tP5HBu
9kxkh9vNR4Xay+t+EhFLUBShq7r0CaC1VVfeH1KLT/nqbsWyCbIglCNyQo9W7UbN
99JZ1X6rsgUfwo0oOYdf0CnLRXh+/gjtG1dXD8CAy0Oz9TXvdY7c7+pA1IDa+1Vh
Ig+yA8h/bP2Z04vrB25DmBCPz/gdh44RwrvPcjzWMcUqSH8+hNs5VspJhWfm2tzV
vEvtyrJPQqjoLpanWieYApLs1pXpJJRiqnZ3jh+SjWjutooQshv9MfeuCDgDq1/t
xgjpe1iLtWIVK3H9fseao4W53HzSYhOjT5FP3RUBdeIQo3Om/54qJGRwoHeYJ4sj
Bu2EWjBc0FevZvAyJGGr7+cqah87X4XoIPTlRD7jJmwmVSuNut5MYhm9t7RTaWq+
ffeVict2CS2tWyYe4yDk7wQVa8Z+7fcGJgvjDvYs2OdyoG7sZCY61Jax0lcHw4Nh
6vyeDV/SV1mgjI4f2Njd/vd+nR6GGrRYsfsrcUqZgv2Yd6HT7kb1VjH471N0UGvy
LF1wu5AL3IEVPMq2YkDXCgdaMdXbV0eaMJUnwDpMEZsKF8x3nyhMEnFPWsrymi0Q
gSwNWVPrLo4STCuIVFSaCsmUL0KFYSkXGa7XHecatQVSZDJyw0XA4i7l2XL0usIg
JhICkqoMltsIEZaknxKqQE1zFyjmP7I0LaUOJP5lpeshvN3Imfeh4TcSwKjYt9vg
S63RRfjWZ6IMhCGBO81MDJtX/7EK58dGNibs6WCI+EjiWtNn1J1xwmpw4fTJ/xra
BAlt84p/SscLtKRqQ6v33jt/ovsap4eeVBrKDRAojMWZ7ZCBsbSvd1rkkqF4AOqL
O3cpptXvan4M3tNZekzCn9/VzIGSy9SleZrfOWE1Q4u0EpoiURHLzyEHxgwdh4bu
494z7JijHSJt/5dRb5i8DSv7yN8LCy6rNiRI4Q0DnRb4IdUz7DDwDGyJG4OdBNRa
3Oj2VsWEwqDuWJVU1X3bzslfq7Gfgnta3xv40rmzC04vCskLSmptTL9/9E2DdyaC
cZNy7ABgnTiSfgIL4JFJK9Ue8jlDcSU3n/sUPtE9pac8+9nv3vJKnAHDOzaEINxe
MnGXjQ85/jVR2q7xo/zgl35SamB0y1+WV4+SJ2x1z6Je0LUjmhXdTMYDQU0Rtom5
WviftbDG174rLABYS3yTae/A6cceme8j4KNShEIvltEPv+66T1YbZChcqyhGDqd0
RhOjtGkAPZkEq7AcHVwJbhc3y4AHZafzcSF9hFc92BHjuDygiH2wbUpLa2bUSCxR
ARHJarc6MGr1n65JgmowmKwFTTxT+cq/MO4AZ6LaMM4dxxJGQ4nC5OdMvTopPH0/
IhEeFdSBqfsW43ateUNSkvHDQA191tfa1Bkk+kr0DrSMwATSG0eNYFgV4cRO4q42
RY2bH4AzwXsX0Fdy1gWsAxHuielLBDrcknA6/UrQLf5tR53DwlUBRcClD0WUTaKp
82nlSlX69Daj218+puEv4D3D2hhfuPlB4T1l55LajNjMyZUm+XKbK4vY83CLg3XP
B1cxDEBRAdNnHneZuGUsxIlw2No22Y78yI6bVGbT0CMxdbZVf9h2OemNP9yCvg4R
hxuj5UkDqsqXVJEl8ZlPocH4J+sGZXPG4K92s5dt/zbhnd6yWsbjuGz2vT+MLbZe
Qb9uxFygDMXxS3oYZTIToPQTnh3qYOCgwVbWSemf6+qwuNn6aXrP+n4FwaWVeAS6
kT1HuiwsEuZbP84UL/DZwcQsDvKZ85+kQTMj+OXeU0sljtXw0Vek0avyKJy4i9c3
DHTKsjY40ax2g8/SGp51cVL4vLrMf3WOS3VZHE+qgAdWuuImYc9nIQQbmFCc1cYo
L0wO17PFREYLINyBJ30imrSh7SksrC+iY4r49M4UQa4M+qnxMv5q6DqeKnyFqttN
BkLlIy2MT3gOZK1rgg/+qJxq1HX63AGaGY+WRl+23zoNh8fbaG3TIYkUbRF68g7R
ypLtpFnESeKbmIiYbMhkL8mwqG7RytItj+GrFkot/I96A9M1XNFa983+/rm5tmeJ
ttnnkM6JBt+eJj14e7uVY73Fp6PomummX3gZaUg6yJI5I0yv/bVPW1muvIK5uCha
gDIOZB35ICtwIUqWKyqkFOCzIiiv84Kk5pPCoFM91+iI+8mmojibGu/KU8ujxVT0
Wrf3skvVgaJT4bzyLC0rRMjt6+C7yo2lwcSk8SbYzYpq9tJ77lBJbBffJeiNH+x6
7OLkY68e3DoUy0Q4xGpO7b1G3YazJVsVjSQcd2kZ7RLKb3X7l5inIEU8PqZwUkW6
ePj6bF9o3ly2o4e72iKja9BtEXvliH4dkdK992AKq6lV/AwIKsZOK9Y+eLrBfeib
1bRCXINlzGz2gfcAjN4AkxtuTeOdIpk9vtqzNtZHbYajsRPftMrFxGIhZ6PQAldS
aP1MIGN5RmrggT6gHjJmIzmcZvTEw39ez3crWoZoXDpheAW7FMGMyJYMzejIEjBu
6kXK3RxReJO45ii8YdgJ/zgTIOl6hEzAxB0oyBCJoVftzA/WdVRyvtM/Lx1flN+3
0kQD5697rztsEY8cuEF+vhMb7oQ+K0b1tPjAU0oMGXTMnJfvtZCLXPXZTikPXOi5
jY+mGrG+kU27w0wh5orYVGjmEmrbyh6LJdFu7vJ6msWsMdnjBdT6bm8L+6lm2ldE
NR5DebQfV/VYfdCtMT8Eoe8RC/gk36LcOYN/sXsEO7w3dI75z/cgxuIfyC12TxyD
wbn+JGYRGwsnb73XpFwYiIypXkX92c2HtjArbvZVDpLLrslkfOHIr82IUtpp1XHD
08jBW8ngpcWtb0SJB/aMjvZu1rGWjcASd7+qOM2lU4DrzRIYaw5XV0oBOe5nAhi0
8KNX3Sh9jS2aYQ5NOQE5DloOZkALUrpBqzOFv4amNQpmWRRlVIyM+0uLmHaoiTsu
TB3dxdjPFVOEcDjwOC+8eMLh8yuOkxEBTAQONOPgIFXGkhd5yS6nSkV0FaZDWsUf
14ee//8L0sMarIWFR1eZirZ7R6DAHKhAVeU/jc1MzjuoIv6tIPIA62GXqzPfySNG
uCNUufiiLMcbh6qqyo+t7b/pOJ8lYQBL69GLqeVx4RwB9gK+KOGBfVmaYP3xlaiE
VZI/aBNXVal1THB7ENxk36rY91k5AOm4l1TRqan0rZwHKphHAwtaX+OTHKf+6MRn
io6dw+8szkYwsxqgxfyOl7tWrk+OUkYZLWzgHd5gcSOHLNaz0jWkqgdpHWhOkIO5
mOLOGkwpMHv2IgkjlG5x5sYwcrOvXMaCiPQN8EsPXPZ9LG33x1j01zfPHgEBOW3O
/OQNViK7sGrC9GkAR37u/wXeyxJ9Qza5NqzYGykUkAHPdn+SN0ZsQg0GI/4fyT1L
lTCmeJj3AroeG5qaI4vDElLrETzUeYUKr3CffCMNm0lNEigfz5003djaBDsN8kBK
doalXyXhW/ASt0pMk9m6UMmf92wqxd2KdkYvcqE104h9Jl/YV6HZLK0nC0Efj2yD
NZGkP3YJrfDBVVESJJzXfvTg/+ch6/Wr6CXxgq4Z0oafZJdyMBOv8GKIckyjZrwF
Wzxlo7RdN0v09eUvK4TCOAx+RsbzDUWru6fHD17YkjU5F76aiwLyBhzkIF6rtE8u
FGZGjlK8GEGvoRf4G0K+fE68nYi+/05d3AnBTH6zpBw2wYQEhVZR2TUXfEe6QjjU
PIVR3L9TOyf0AuY5/3mVC80wM8Qac3FMgMJzosAjVSHneeDQg3/tRh1j30zBByI2
Zm8yq4QxPaAI7SGF1UAfRO/0UhB8dM0BLwZiHfrnVqjkdJQRK95FmcA/VkR2SUTz
8d1wvkxbp/ctrCFu5XEz4031BIZDcZS+CssaRmXBmOmXQqn1awTXskP9zqZLcc13
fxlV4ODFowBIJCVPyjsWyvycAAp9DqHYLUNxBGw2q18PLnTmJGFmDNU7yhger3tM
Ghtcr7kvI/Ne0war35KbRXvPDQ/w3TAHX92Ln9COhEKCHLtOx3MHv2jSvZS4+9gu
xL1MSv/fr9LC8pQ2q2o09QZKx+BwBZIkBpASo0r5oqc9VJG3HuFVbjRMdNvWp6Hu
rHI0/L0rqzmP2z6foRIEthKGm0/IausQGV+KxL44WGgIJSycdp53vAbxZRdMC+7v
uBXE2/podbVdvo87FxHXnPR3tNFs7prGBn8qVz34UA15HtD92i8gkoYcw94X5u88
SpBQ7n803IJIuhlsqMElYtAcqmDLaQT+UdLIQUsL8vxiCXinvGDc1ocwf7UuAbFn
TXYSKqYD77RDRkZ5IvvNsVJ0GAXsUr1d9XguRjONWyogs6aAegYTWp7XJwnq/1HD
vMZ/HjjO+gMBpd5/Bwf1IlRUTVDt4j11U/EYXmPraobA8TPxN75mDv1gH0YcKI/+
phlZJNQSCsRdb4NSQcNxS7ZyaOEHgyNvs9P16kNJ7aC6LV4vuDzPbovX05z5kE53
eK3FWuej25B0fu5dXzkZ/rWBeSjzPNmA48jxAZKJhmbQNm+0pJmT99lWI7+W0wtc
FMLqCqPD47EtMAHbN3Vly4zs7W7Be7yX66to7VN1j5gG9+V3BTNUoo50UxQBx10P
tw1VUIAb3DoSROOI5UVToWSwJUsCnnKxIFHV9R4V/vgYlT8Ff3J720yt+D54HYzn
SXTQCMHqOVI8YMRuaKR9Ou8zubQBO0qmysA08+N7rTrbH4IK8RYm3D5AMl40I57x
aDjCA4ZneOyFp+kb+JpdjAmOn96AkitT/SaHzuNgHz0OwG6e+8n5x4IMAKmId032
I1X7qcA0FMPbTgzkCQB6S2mLvlRXzV/KS55DrpNfuVkg461eHtzDqMOfSfx/BnDA
ye+WUpV8sNLd3eHRgdk7NEPBOQ+LOEsBH7HJI+FLAr2AckoYFxKO4TrXxTkDOL5N
XBpB69U2yXS92eTErrui1neY/gTQ7UcLO5xnkkZfM+BXjyRQRCI/nddDqdvJVZ+I
JKT3a3QUgKP/DNZLt/6QcEzo+29ZAdBZk4ZPmtz3lU4ghllJ3I5p5EB39Rh75Z3e
kCK4bBX3Hrq57padPBj6Vp3GnnGAe/4CG9YeGc0ZjfAKWUwbsqKa8e4tZbmpilLM
xV1WLr6ARYTjN3Z2wHAv3PxNk4lxZC+TUt9yBWVwaLE70chy7Acp58D3kWEtoZH+
+6QwZbPHKdCHLotDG/xIHY7JB0cLqUTuN8wRETs1aX656jL62l6a7z0Qz9clM0Va
3d5NZoqZODO1ykQ/e04hMmFhln6JtbIDe3boUuvgM19ureMwx/KJSss4hXRWNGVO
8x98f7mHINxlGQ4EmIpzfJZ81iwpdTOzRtsIwmAfmYvBc4Es+iwx+orVTt9DAYUw
H2t4j8zS20+Q47ixABgdTF4a+Iq7Qzg0uVeCGxvlMpS2Rx8KHvNFj9vI6/9jsqvs
o4TO52a+jnBb6BQJ0ySJj8/jAA+YxauKfhGSX+Oz8onbcBexR06FqSdOYooQdznt
RAYgL45+yOZNhoDTpDS3wDayo5LLviQ7XI7kYs/L2Qd+ZXCWlL7s1hB/Gj3MOmYz
JYDJlqK5JdsJQZztvngFCm9B0Z1Ri7rpp8R9wzfj68KD9Uz+1PxTMOxhX/VkUy3U
M9Hf9/nIc2Jw6aukcMV/Imx/xj7A7GObf08ePgu5h77mYtiJ7fvmO9gW4UPX7pbB
E1vZW/N1qSE0cZAg6KBEnzDMqTKcvRqgoEwVsvAeGPqo60zveR5TNrk1NIbgYkpH
FHyt1ab3BS3gnmUuBp1X/dzie7u2h8L5WDgozOft0gv06iWqIfTdAwY9q9WixQYZ
0CLAPdaficEkIWxxT1P9I5Mtp73DAUjM7kOHY5FsqJ5R+xI+BhWW6GRYMT4VpJwY
3YgbuDVxMQnZ5e+EuTeXZHrE1GMnMP/I3MYRE4uajtMJDgAQENSXz6ymhof945GW
io0Haq1VgMGuwEizoIi36JWCCRX+0yvEGDYDYFs/AXQGsotey4iJQx5bxn9TobBX
AE6gpvaCcL4yxkd1qEjoFzyWFZa5K9+QEPUXsguw+E9iBrcbkXEl4Z7SAm6zATi7
BCRuRkg8LA6Ijl2uaR23gRhJexzXfrnlu4n9TWEa3m7zB8Y9x9xflDLiqL4pVrTr
4J2qOeCoY7ZfOKLgYCH310vrIfxyy1SzvvLSGW8aBxQjt8XG70VsjS5VmvOmb15x
YJyg1jnYdJxad6pCtrCNvD2RtaZLMlQ4A047+w0zHfqEc3sJl/gBZnwN1QqL9jVX
K+gf07C2NFtGIQxS2ymBGEKWOf4O5eSwneUTPiRIEQ7UKJU5oYWPj49JgHaOeFBm
yQYe9qwCI1DkP5CyqdttAmn7PaEC1AeVnm31aK9oLxjQAY9v6HmMXXvT5OOybS4p
pWu234809Jutp3WbgHRXX8lrcfBS0F6EoVjPlTNWLz6mm3B1qKXpjNSMiAY7MWCo
OjsKSFufyuNoeliKCrhV4ZoOVbk3k5pu7mYT89NauShgEKC6L5XySqv80CRd8uwK
sL0LQIontPRU8XURPsw2JkSEezs+RhvjAyWaqDqWc6U64wJ5EnrWMNKN8jCv0egr
yACQy3N79/yl/M9IvBIGyCfsxtzEn+/MejCotulGWA43VKkq117WpaxkZbYNZc4r
+1VFC07bbhDZUDEyiinbvvDaTtNyGpVJBm4yxvywB5c3UFuW3GWYG6LQ8ru1NeWf
a/+jdjqRlb8gSDB++eRS4BqAiv4mb3KpKbZCGGCg5V4nF10AIwj9Vs6E/u5eFZ8m
tsLUc8BRROTkE4ZLgtjIgYoW+6mUlF0QKSLUuHV5krw2g0619IP8fA2SRbzDEp7r
2GDg+l2IxPixoihCVMKhA+rYklrstbxzmqvPcSJVloGASxBRMZKezROdvpB6QoeI
8Zd+x6HbBGab6zYUf6XNyKARF+z+OLYMcInz3FLmUYpE8Q7xMdGl0UEzsPazN5nA
ezZAwF2JCLsMKNacJg5Ffrr8C07r/8vHQ+lK3KX7bPvQdvaFDjhnIGzKtAmvoDp4
qb5SBFVKdhIJOukLpGkRTE+Drp3E60PnkTMj29zY0gw/nii78dwp3uBQ48UYjiYZ
MLfgq6boTvflVkX91UU11rTM8fAsxyliKE7p7IfNh+TSfjNJdKFasVxeosqARUuC
UNWCiVDCQrPW1LHgKIoO7i8k3zx+gZzYGIPON1gV2+qaxMt67UqrTGnCsCiLXlTB
D4lcqhmyr2d6nNBJRsBNeuwMpfbBAtFQsx0tzKrnoo4O6sg5lgpsbyTXCOXcCXkz
cuw5rgSISJXCrw69n1FvlSiSW4Kejrp5vYI8Ilr0AEcvBTvgabj0aJgFV+DTQh9g
F+G7Z+vVKHHtdfLoSlZhC9xOwX9EoHUnzfcgHc9MoxSFF5xLEpHFCbtdfwGwAGix
tW44UrdPBSBTTFOBVkxf299CCAMl+8FaMLLFqyOrqU7CmffGPN7iQnyJfxaibOJ1
bsWBu32RZb4xSVUzVroz5NS+yBLqfuARNIk5XxBctm+yLGQtqBS/P/29VsgK8h9/
qcQEQqgos75lr2ZgnWCMtPZUd+HjuCpKaB0cyQVo4DVH4CbRt3xtetXKrvHACR9C
1vNATltPaG0YT8k9+GyIRQ7Xx2etdfCyBRguAbdHiFwPCKFovWYlqwD4Nm7c/X1t
BGmc5AEIq09GpkklGRzkrwkR9xGy1JrolL04gOY65unu56aY1Yw6sTm8nnf3NuTV
HMwj01pJOOj9+IXK/JR1VzTcpEvfauxhCISkuk8KDX80aHQgs3qORakK6+VPpFWh
FIFf42f88tSfdsgW2GMvpvjnifkvwF9gIvLzD86uMI43sbuEkz3TtUAASQ6UeWLN
j9HjDl/eXM4x160+844y/klFvFrTjwj4y/bDuxPhQOQLrmR7e4RmDV8mHHZI6gW5
JPrg4hhoHm2IwyA6nU5KFii9pVhmZadn9g++0wyqmFg4OFvnxI4QaV3gJXMoRX5y
Dy+DEwPgiudWcnh0Cv+QQaU3UwUBm5jIJRbivtWaWPLv7mgnk705xURvkgfC9QHu
BFy6/S/0HQkLR6TkhjwJ2OtTqTuooRTfLoD/Ndthg0RI0xkE8Kgy0y9Hg7HpGTMu
WezTTOPP57TIdP+bblShgB7qCX1ydVYqvrmgGRu/zsHuaYa9ikVu5hq6WMv4Xc1/
AlW9X+LKL8Ess8x1iDkmoyezjtxGarJBhD7DqL6IQgnQq3C3oVEOglhKRNjPyJZv
SpjEaTHUaagU21PWPs8+/MQycVswWBDkULXgcBkDOYC65F8oFPYjNddEOWK7ArYL
rHPGx+5rJGJa96RrMgfXDErev4MP5Xx1ivXRfLuyTKSBeSWPGGSGYcBDdy6NIJMx
+ZV/Yax78C4duQlpMAo46Owk2JG/Q0rtxFx0pqzGhgvwmnxPfjmE+cP6DhuQzxVP
2Qa7BJUEUYt17nZ8BgIXYpomgkqZeIBX+FSGICrHOLp1ksSmM2Psy5X1N0sxp8Qw
SxKKTvfbbSwLI0oFcROxl2AMHbFRV+lJtEnlE+odaQ2t9MgmL3Uw2IZ/dSNIxF3N
ryLodS5rCkQ69LX+U17GDA3JCE2Q5UywFrksPCqb576lDMtQ3y4p1ueHkKe70GmQ
ezmZDOoIxmrWGv13Yq9HXlCz+2Y0cQcM98YWbvkxV/V1ondCa5Y9uLkLcTms4LqF
Jfyu9IN5joaXHGr9VsvXluQNy1oluY2S+oB1c0NNWdk=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bUoQFUwIHct3u2KutMv8ecZfUv9QRCrNupNvCa0mbU34/ukJqCNy/LPI1P8gC1/3
0JnqH9s9Z5WYInhm85Y8R6akyIDrrfZtJJryMD9FES4gu57jTP4yDP0c6udyiFuK
25hVCFPZNhsY06klkk4w1+F6jU05qaYQPbKvaOzWap430HAJgnzH90OQIkL4+Hi7
AL2+lzSG+szwCuYrUVVTcbzwNJvjTixmGBZnCIq2ERiO4/UQzqIze1vucM4JRyqx
2jlzNJwPvMddY9yvIYAUIC4eOg75H0sV2kFXO4jKnM5Uy3BS+QwV1wC68ijVXmNj
9qQ6pISn9vuFB+WL9rQuOA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8800 )
`pragma protect data_block
WZBrfSLUMx5LbPHblwrLbklhG/ddd/N0+0AM0xgUN1o+UQ11knPNlpcOR7SNxRvg
MdnKBumkVx5p/MHxt7LzKHMClVOm1aYZcCqtWhqmrTENUi/85I0URS3sxlrlV7LD
oiNvkO/MwKtc0dDP3OcVFAsEcgELahHq1sL7l+XWOzmRhLnAtT/etKVU1fLiuIm9
Jt1FflQc3KhVXJfdcgjO3Hx99Kx+jko965I0+laqqcuWmsmYJDsPVRC3E8aIdpUF
TLDtdFiZncZbfq0m4DM8Na7GAfw6x02bi8d+17Mx9Xev75D/mZM7uS9C5Dopc7Rh
rK1MxXbuS+qgCH8HVmsgbSQWXTuJW9WAcJ46AJmZhk9O6TzzcwKYvkf2A7AzfZTH
hETkoUEvN7a58XGAYdpf97JVjWQKcxmMVYkw12JDpd7uU6pjR7uTnQPifVCu1fb0
+CFSPMal4R86V0W7cXUvKsDRrsZjn+pyAiidEQ5qq7LSxGaI+3xDCoPV4G8Sx56T
wgaCwIzG1CvtlKdTZw34SS7+SAOMb6j4VoyEolT4wPQq8Gpak0De6KeKd+zilvPi
W1+E0c+iL+Fyzzh3G6GWQgn78kPzgLCk8vmyAXTn/6gj+qCs16DGZaksnc6TL8jX
dW2uo7R2YN3n6mpZBQivHY/U8UF4ufcgW/uHlp/t8UcEJkcT6tBbifCqrSZgqWlO
PckqbZEzss0VYk2YrmvKU1xyrFfZUFvQgaF1Nq+zU0XZMDHHJlcK/6+A99UY413j
hbOJdhnkDHPELQV/W6qb4NQLfMnFKjkBRX0CLxH0/IpG5LBDvLg2/kj+AHqSx2zU
GGkW5OHQuqBMlVHSztiyN7yVioCAgvlikrq5YEyBW3/kIRonxjjOjK4B6rsNAEtk
/HG+0WnhgcEjyz+RjN/mJ3sjnZOGtz+Km2t0c6PqS39WnF8mm1FlMaKtauaNH8Fx
I9XAK3Dr59LJZW5Fk4oYrEowYRrbyIy3lulH3X/CIqapjouwcf5PrdOTSzxQdbhK
2ZmPAyRdM/O0/rYG40AYp+yzCdzeLcXqKajPjEFDGCLF268Nh3rguJjeb/jJqA3g
dY0ALwAz2qeTWvIsthNhE2ExUwykCcyQSYEq0Wqmp+sA9u6+DIUw3XBcq8tAqhgP
pF2vA87el4pVAiV0283LqCIFhKnroODbJXFVtpgV+d/Xg+L+QSvPrSLWY6qpCBD2
45lhXRBcyOiqICIxoe+N+pc8vETcbRrDPdsFYFkCXjm2zQpRHYapqV4xjvuUsa54
dp5qOOlZrNOkBCBzTSA1N73yd3xZq7vH6huSbtpWqM/6/WiiI2L7C5Ssij8D9uzq
DnDYNNTHX/vGYBUNHqKOnjk2vfKopYB18mXbnSdelFXsMAAyJ4S2+STdziS/dJcO
XjLW+xzvSFeThwF1ftlo8WqT7++0ruXhl3FdXhHhJBr8FKoRWvt/1WaCAqYqz3py
rEqbTc9OqdqG8vAa5twP85ICpWle7dKmONYHh1Rr5M2wlAngC4w4wuSPGjH/np5G
a4V6JibZuUdbiGR56shWdRH6rf8QE5Af9QAuXh86B27wm0MlqJv/0MO862KDFVvx
jkd/oWr0+KGc1+9w8vOunR0+RIT5+L4dcKvLzpFk1jUiNn4uMSzB2t/F4BEtzyrU
XdETx9uuSguXCRsWZlYVhHMeH8e+HBuKWHvd3WmKZf6nhXhLrbhXXk+PpI6QEjWd
tBw6j+C7RXEUsp+fDCJ18P36TC4axucTowsdsM355U8mM5ESnQfMF+KYiCsIPZI3
jWdB7KRxP2FHahdk6bJU8K9aMfWjixyf1ly/dTKj743gio7okXSfCz7/ATkcqaE2
Jf+W4fFhy25tR7H55g/4MoK3VpPC1xibI65TarccgsQgp09mc/+KgYdZwCZJT/ku
QJoHMcXiRGB9fMSsGvkOmy26o9zQ6Hkb61B7TVf33n10l5ORjH6X51Dns/RwOvl3
GImZf7x+/1gbcxCWAUP4SO0UzLwhGapisfb64I4Z9gacEmj4US6qdTptW7aLG0pP
L5CVmEY0WIIGzjTaNk5X4tJrM5dJSa6gOAnOvdckICJMKzXos1zA90YmPXfCg+A2
m9XGN6NBCgjYYBYNj/IwizNoiNj6dXdG31VXYcxkXCH2VB3PwCdtMkueeNYNbrZ6
KZD9y7gpP3kuPc+sRStc9SBI39fG4zhKQL0X3u5v5hUUckP6RIEvckDRI8Y5eMSr
OHO/NvBswJxrjgm6U1utcePkdGXb9OmZYtg8UQZQZgWODqH0uNtkzb5IgBcCONu3
L3uZpbpjLEwTMlj5MBCuac0G13FGua1FVfbt2OavnNDXI7VtMqSJBnpm6E8bM3ne
XAJl4dowHv2elIhFRTS/fVaHtPHJWOxC+Es0ggHlOAYsJOF48mbRyO0Cp8hKoxjC
2RRaVg8kBosH1KAOieCd4D4B0bM7jEWEzCx0SctEIxAv/dxZMy9dbbH5By9uRnqs
BJtGXs9QTNrHtS3W05CRnKIbICk83Agz+xnAKTIpZ+FpVKHJVsK81gpcfOhzIvqA
ChM9resXnlX5cZL8dAa+fQ7TQs9XREYPRF66006byB/dFJI0ufSv4/xMW5iTgccJ
4PwZBJ5I+JFztVPHmIQOVtDIGrt4goTJEqZd+Lozzii+BXhylpI07xUzm6Ga7Hap
TI8GDhn3f3+94XmIRFyO9JkZGxVbvZEDpg+I6h3igwoDOmmteM+6eAgbpSvREyyZ
fDHs1kE37DwRi12GaKxxDcpWW4HK87vF5lit1M+jvxt71qwRAFssozvTO9Ukj3Xi
3b7EcNiGdXXSkKa0VC/AH4Iyc3RT23Av14tRREGh4oC34pL4p5vfEwCuyDs0DlQ/
UX53+goKK/tSJh321/KAyqfmsQ6ABQBPxOZzMOQXkqXOdGseoTb8N/S+L0axF/ZY
52ell4gemj8Q6WHWT3sBAaw7613YLUimdRYUblt7qA4+7303BUogHK0Pb62JaZZc
FWEJpSp7UHAhiTYMHA7wJVPCCQwuPACrb23M5VfUhHzjW+022oA5NavLg1n7iT7S
ZiLHqqHHUrwr6/mBzirbO+2Ob52AVAEeRDDwSSIAtoi3J+tiOGfyDRyMXes7usFz
TsGJrrMAx2EVQ/9Zx/vCt/WaDZWbgXKw7HH1kxV8FY4d5QiIr7kkVM072IF62xuE
K9aiAmYkmrMepyQFOBXc5M62e+/ZET8TVOHr3YGETCWiJuC3XGWF1QxPbiafPfLO
AdiHkENPdJI2VEquNoHbWDuWDOqb1pMj6yWHyAEHj8MQPBc/SMwEDwNlbZ5Ti9T6
RvL1HSkvGP/4+pOSM6LD/mJ7RG6z65zq9no4ULH2mSSD3N3p/O4jqX7TRB7mxS3g
7qXzW/e5JK6BcQMg8ae2Kl8THH6MvWI94ptcwTgCcwMl/O7AZKMg4YJ5dqFcQeYj
zDVc8gaYUoH/UEjI57TehNc8grjwQOmfSt1y31bYU9vXuxeyaRuHNN6QSIqPGgwj
NPpZXp3IGiwK9n7z/3OExtKbUPMcptrQsAIcQAGUz+XPzTdYGq4R5QWD29g5x36I
V+jlUgXp2M64LcNzZOubNRU6dQV/CVwHRuaunKdWRmvWM6WxOsNRxNo1LMsOW03k
AEEvOcefNTT2YV2PEitbOElhE+z9GkvdTC11VAu95xeyWaEimC9CgMWEot8EATyW
N+rsZ6+kikt/GRk1jw65Lmj21PJVqxKlUIdL4yQAKk9Hjilp/F6PWXhlmy0/ufKk
wfDKNcpkbK1OOwUjgyojH51mUlqIN7TcmfIqmOdSwUgnoP/5MQCYxED6Lbq/59p0
bCtR21IQICXuC1qgbQaCJ1u5OOEH9jzcMxCrcmz0LO4o6dJAeAa5FFm/rpwBjp7s
q1UQQaHtsyrjYMaeDLC1ngUJtPBpIBgjlAGvPyu/B/G3S5vcKcn+vh0VZwT29umU
RSLO/gw/BpabwBuqW/AfXCCMqxXTpxyJ+CE/EXiVQbQie/rJ9uvWWbNLaC3eznVM
UDETeULxf0+vn8gRd3S25uYY25mX4sV0ssjikVQBXEYHMBkYn0fKoBvE13tVQMiZ
S8OQ0ySbOt2ywfRJEID6XznRnXH1u6rbMkORr74CceKei5e44OyDsxVllYtNa+bH
gQBWN41ksR+g8GKQW+PT8EbCOmNm8vaMvv04QXZDPFCsSWBfk4uUG1cULIsBeEDn
EoFjlYRm9EKmHz2jxuet8JbcHBsJPk1MQD+FtKhg9TFEH0ucIVNpKuxnDC4SWfTB
tkPvdxdF0dalmcgQO9GL3ObL/iyqaEKet/Ywi+gJTYpafpqdi79JGOMJmr7CsHZO
3n+wdNCcbrRGytt918ArwdKmbKsbdYDMdiw//IizazKClQBKaqnyNz1BNV5fdKcq
EX3g0fRYM/6xVeSwG6CwIV5QB1hJz9DOEiBZX2quzPXLFum11k7Cd2a04FMTYC6J
SGfD7L5erhOmIi3J7jo9uy+b87gi3HcPacPQfKXuUjOBikJX2r8sJ+rhjEnhfnVj
AiLrI4dQaxqsT4yDffSnQyDvcPRlboDWLS1mtjzAfc/9/33Mg7+sZ2mInQo2zqRU
LEWwzm7QjpKTix3hk56wCRQExU2L1hhwzRa0Mr5ZPKbu4nyWktLdudQ8vLnx31AG
M4Otv54HITDgFiV1zTuKel7Vzy30FDVzXVbYjp9pbPV8PYBLcl1gSw5Zd08SB24K
L2QjOalpXMO0P8aG7OdhugkpSh6Q20cjF6aJdnpA9s9tPWgjKMnd6QRfDMRPqyCO
CmCu+ns+sgiCbUKDJBukLAsJjq+oQc13y+QNwkT8vS4dku1OUFDogJA1s5ek8ikb
zTE2cd9YWpMHdq46QpI1dl3uK/rPMnhGUTOE+eVJfta0iN8/lt335WcR2qhUT7Kf
4imp/zzBTC+JLrI8AaSBaKWdQLkHsBcfXLmcXg7EEVslYHeUmlWN4aLMZLHLNZM6
+3OZfZA6Df/mm46ElLu5uTZ71dJ+e6bmtehD7j/gmnkWnSty1OTIdCOCgRET8vfI
DS7pE0Fd3gkn3XZwzXOzbRf2twiUAJk7IPMW4SX7Cu20SkpCFIJtnzfBkXL3umc9
3tFPqOM74aEMfSsc9RkiLYAvbSOGHHrNdWKfqIGMIxzBtpVsMmAW9Cv2Kfv10MBa
zB6LKunEIKQFinaI5sbZN+YHsBpaxds+LCPTasihLcU86P0lIh6JNkqylhQCdsq6
Fd/IBJX0f4+lC6X1rM5l0O/hyMpWbG4NqzMbql6BIxRjKagHFkVcFE6mse69TYFz
K0CWRtxTnraQyUP3jQndKpal8eTR6yn3R1H6Xlct+9LEw1GINx/rS0B3B/W7wdeL
/z5VkmSlGs3HwgqErkc2Gl6SR3nP8xGMm59t4IszyRrWXsKAAgrF2k+ne6uG2rMg
5+zI+5H2cjxd/hIYB9WQrzTz1NPINj85bQUcxOPQcwqoyDze3EMS56ktyQmMoJuq
W0p1p+yIPv2hkxvDB5xK4nmtre5BElJcJ1f6ed2IZUH3L7CnJU713xNg+8iXvQHG
mQfNd2GCd0dWzMQ+4rlbCnZyDfb9f8oNijcDUgJLZ59Kofkn2J72Bn2ZDGeuQldy
FzvNJ9XtJLuwqTLnw1eNZj/2kmEUmachLcZZHzfCKFdRDhEVTF3O3qBanU2vE/Ma
2X6cy44ZST49F15CUWK4wjm36whXdm2i5puJ3Ly9HdMLSeoEeXRQg5aCBj/XRwEL
lBpaNKyVjqjjKSNK+idHcnrsKxjPhIb0gfYIBo6yL5qwNT2HoAUBd8vL0zvsF2li
sSX2Pxm8gzJFQewbP3JZVH15k8lArO5go6YOMw6YBGbNSQiBZQDKL01B6Xxgl54Y
N3YJNV72AjQNugoAZJ0EXhjDBdsziKSUBPUIXxtE6HYMwCVh2TepIllM+4x7rjt0
IQ2qexLWspe2Tg4GgKx4vZHROE6HZuVWc8JAD2IGwE/C+IkBLTSSQs4nBkcJ3zZG
3QI/J+9WLI/M98ROn8F53/magt7JOvFNG0xC+SLbdqu1VN957phSO1FKgp8pddTh
pYUFMIMRFNfzgI0eRyTdYdYkkmTMF5bRb03DMz3wwB7pyHXYw2NCjzgqBCm/0X1E
N4TRatrpCBhaQuWLoc7rbNsUztz8d1ti3sOH5uxutoenOiWPBLpwI7vBUKmG0q/t
wG/1VK5C2hrLxuPW58gY26iXpluasQg0KLSs6g3J5TBPmdnJyf1CboZb6d2POD3B
VTqfYpIpUYNaofHUjVH8jNMltS2H3tOg/akTCUloPqX3IjZersnI4NZUKVNl9ZHy
0Msb7VDAvO7/5RMmwAPV02/6KTM1oCNwloJ1mWIRI5ASF2C2FhUgwqpIhXAEq01Y
UBcYMD4qJyPXlHQcMCka7uGlcx7yzaN7tb49pHhRGTbBOSkTmvDHXaDdarVE/pMJ
SMz3cts51oMgRjqVnjuNx12N19WA1QJRMScWEXY5XEo4MtvrokJkSb412wnOJnRj
pyWEffFQ3LMp2kYlksp3iGv0HS77xj9TvbdA+CBrb16BIyL3RPjtpNFvVGsArTl/
yCJRoKqE/CW3hIydmXWspRTLitMFwGT6k4f7SQbkrocK7+5ityRVtDgkWd14+Ouj
ldhdKqRPpGxXgYBPNiZranzhJ90YR1hpd9rTtVcBTtG41unV8aFHDU8STRecsYS2
VAII3oafJcGo2fXwd9niIxCvazSIoOx3qwJrRsiOvsnLNy2pYn2xk3gwCUH7Z+Db
dOzxnZMHhBmBggc7zHuFQzlaAMgpG1+oHdjgtACu+xQSZRsnVMswv/DrIGpX5QHH
+Tr+mCAwHxkZogW8HtEAuYE9OdrJA9GfhmxEYQOePsNpn8MOYlD/R0It2tiJ1mKO
vUTFtZ6XvanUq7LMV4ZcCmg4UjSgXkvkIyZWQENbqdLgDmaiuqNl3uLHBHJedDVm
e6tYz06pfzSEl3THZ0YkGFY/4dD+UK0i+GNV6B8OGSCXVgcZVzx37EJBQefFU4m4
Qnl98fuc7Uk7mrxOzjjXTiochJEAvEdn60FTpJH0095KUO3E6GReff5tKwS3hf4f
CHWgOkrVpFOPG0SdCjQ3C2VhHdimU5HmXjL3j7K702cyHLPAqWQcxxETR/eObCic
dWMs1RJLkyyb90m08hcvxReEr+MyKn1tzuuC1GcQv4Z2odNU2qkWPwvQz26RMseA
k+QobodKAnZIXLMumvLqq//sEaNHeyJg0ppFhlq3TSeQqVr7tTJ9mHiDE1vXuFf7
N1OGttivGJrS3m35P073RsMVyZMQGQIsdUtPoE+9IzAY8UuAn7cIRFNyJVoh1BzO
oHi5nK8sNix9SFuGg8P+ix9mWDKxY0furIrwp6ypVKwk+XjFPZS+uRXl74rHRT/W
dGghFkOBavrBZFdob7iF49WCGG+2JWzAuUIZhk7/JkZvIOARaNi9TP8OjdZQMtLE
OnoiMwgtu3wwIsiNfreyuefAWpJyBatJtj7tlhCcrde6ZU3G/8iQ2BN28l0KrRR8
tTSgHrRcU9uNkZmykOtgRcE+iRWibjq/XZYjglvzVj2ZFMYkeRcnEKcm6LOP/VEd
xI8LYwZmTEaq7C/upYe/qZjMmRxQ+vHcfwyxIzZkPL6+l1s3LWJH7cRwk3zaax5i
iB7JzzYFPAosVRqQkqBVtSMrxtSs2E7F3rzaUQLrjr15G6MtwcMLmYa0KWnTXVZ7
Em7tbMcUK2tyFRZlAXGCdMU7uR7cRyd+ghJXvErBGurViyS8xe4KG5biLUp5qZy/
3Uzh4iIBC8KU5cCFB8dfSVg5fdzayb/20NUp3o9S8agFocEG4yzlzx2AOzNaCPK3
UUwoVC4GthY/BsuDczLsD5R2fOEabz2vdpBpEtsZ+6qkVKLFUMtn1c0lPbN3098M
tJuPyv7fhz+y+ZP4O3okxdQO1XWN8OfoY8aYKSfRlEOx7rzWJzB9FDvWtx00scj6
eBIBDYLjBFjZTOz1QwHUyj6x9LGWWpqWpOpo8TJjKliOpRuKPe1+udxg5SzVjkxe
5DoKz5+jQPzVRpW624C8OdLoAbDn1TAMoo0obI15Yg9JMErbB5yMgMIn6CAWaG9N
Ki64QnYH+xjn+Mljio+pZTPYUFWMJyL6bNYvpO2hOwXkk3reWSq0PSwMyTqGB3RT
gptFbUnl/NCln24c2AH1EBYA/SHzLLNroaeMHYRxJQke4HqUJfMZNQVovDubYrYs
8bedjrhzYfnl8sOsMgcUjq7/uVJLwtU7gIH0Kox7vI8CLg+hNE0QxH5uz227BYtA
bpkys3ivm2j/uiYFsPK/Lofo+iGOgVnx3mH8gsOJC6WX6YFfyzgjPahzufPL+4eV
qPxkojEKyNA2RDw3VWTcFlN9VRuvFeQphTz9eh+z23BhkJuog+F6YBSnaMKm2exv
EJqW4cXrZo1h/FFCv2nxAPkJosLEDTqddczxyIwih8d3q20qS3oEQiCK7gOMjPRv
RYDwC8TN98PDXapVG2rl0WqG0XWBVJi3H3ikZzhdonYAcAHq0DqGUP4LcDYKi7DR
cXRaxNVYDmyAxRgb/78sVRMAJZrU0/v7CCiOO7J5Y4F0+QKNiNq2RhZH9/xLgLSu
piFpf2SPBu9ytI1NWJKzW78mWAM78TSfGfgi5wnxe36YA0o9bD74n2+CsxcXpxoh
fqoGYWfKLuyosiBoalF1ydeJGG3hV4BYaB9kPYn2LZqpISmKLXZPGfEr2USgnsOY
w3gV1oE4Y1rR2nuE5jnL/iFIWB8cyd7itxnktnwoRoLOJVwDx1nwIIgFAY/u7qLY
Jw5VDt/W42FQZzBnv1ttCITKWWniBCA9k2WyMxHJXl7MRuU/rtq2zmVSHATWtxBU
JHszoQaFAm4d4im1bmkaMsBwQiVolyxV6Kocb16pgpTfKHRwuHzoow/d3GsZvw3q
ZHWj48Q2naeOK6IL2283ycbBisPjsEIw1pT2xu794Dp6DLeyUbb6t0RUeNVCtg5M
GlIGk4BCn0+Upu9kMsBN+CRup61SVv/zfVE0mSb+qM541cNTa2pbZPMxiRdCkzFB
0kHeskpsPqrgyEVLgps42tlfJzGvN92ZM8sTBjIW5NvZf7sThiziV+xHVY80B/cg
TlGHXO3CYX9HCJOXFRsQkwkivOsXLZfHu0KA0wbtXktzZYaoWBe2QUW4JLdbHuSL
WZCNOO+KLttIiR5NrwMxsZZAfG0mX3qiolCUrdNg0H+pLu5uG8P7JQavnXXIg1vK
c7HJjfPQotNGj5NSDpTKk56ejT6raKUtUly4Q0C2g1AQXIyGQVtaJGaNv4WWZCqv
WwlhMmDIDdSTqUkBGQDyiVpvaYc22Ge6xjWnkimIxM3Qo2V9q+GYAhpKXsNJ08Sk
fy4xRW5BZbxU27tXDerKJy2r0KLGp1ln+LI3YCwGNI6bADWhEJunQVyuKauVLygJ
ihj3G4iAoehw9L2eH9V9tixPNapxJbUBYVfvwzXQl5UKQqqhtD6VomMkwTWo//G0
c7prfFmsLmLHRnheKybrYqvL43vELfjtBFg7TNHi64GL4vF5PoNSngSMjlu2KdDb
N1JrZQmxe61t6CPp7OycB1QOS6tOUPGyxs/nFt1AN58ulrs/zI19VkBMM/BKN3ST
bLILyE3dkRrhGFuNVWYyYvlXYBhZFdRxjxDFZIjW8dzGbXs3dWIVgE4Gk73l9CND
uxqrphIKjqZ6VcdcS2dBnQxgIy5wYkLihCxqDaNdspv7uksd5PmO8PSjn+HqEiDJ
XtoesAHq6BVwLmiLl3kSzmU5sT2lC0pvsizgsMJYkTgyrokcicSU9BQbNsJFdfLY
e1mYaAsNUP+23/WBtPRGB+MpI4gcbt9dnVEB9678NSyrF3tQhX85NMazOYZlfXTF
w+sfsydq9CCZXSuOe3H8NQeAqlGbVCU3SfU7brtvbNUVQ7fJ73jGY8KF9i0Cx8Gh
Dd08qpd3zLlKr/GgcWnFKtFxLKtCpP4epFnTOBd5005ZOjHLO01uQicKtF5s4eKm
I1jYL9eVT/SPlSAJ3d7cLWiLFpJiLIncHfF15/7wHas0NIku1M3pfSINoPwNzThz
prn8bjMLGp1ZHpYPvTgDlsGdSrvooRZoyMLlh/uays3qUR1Tv4PA5sG+dvIjHwP0
3pkFXJe6+dNP4ENbDIjYenJUMnWMlCqVJcIhEZeQAvcMrHupf7jnrplWc0G1ojRC
7A1DxlzLqOj4VyK40RXl56jSwzq9OoFShlQkA9d9q/LnwbfdD93h2Qx8S9OiZXbp
G6ZZs59l1cRj11hJt30qhKZrPrWINuCdGSqqvetILmuQ31OyTRYlclrZWpEIio+Z
54jh7v9Y/A4AcLkFOK5GE5eIVWEnaGbjU1sIfuMLhlUcL0w2dBfwDMWMvvuTgs6W
GZruBBsnoaeKtkuCOZVl+4SkmHIvQroSNS3WFTq9ul3pKKHTEp1yz5RY8f8oTtpv
YssLBKhRd9doxfvw7tsOgnLKLM+CYcSepocOweHYM3XU6Pw8j9P/jsqkN0RvU7v2
zhEbPSVccVLoPsn/tU0sP5Dwr8Ri43O34dttn/y1HDKY0LuHQttTmCwh4AjCJ/b/
isAWpWhIjZb63Jpp5hqldKRUDpyHfIiMjpba42FR8gCt5/7s2SKAaCfAhZu0YmNL
B2i3TCeXlZlOjsXlZObN/FQo5Mi/jCM83mCah68P0L79RwHhKLT4HZ6uQgQjVYVF
760HAgl2VTKPSTXWsam5U9/6ZUhTT1hgeCPTMWfv8pVbYaDs1hU3R+o4eNP2NxFk
LIgiUNZVFK6qWH3CACdbN27jKSorF9BM/vJ03C303OULVVcaThsy48/Qyt4cYJ2V
6v8QoHOXSfBtLmnXT31ataL2e+7h5NzG2a7/Wm8SgVo+tbbKZJ1d8svQnUbkSg+4
+p5sUknqN0M/3c1h8iVWdr5E3OStNEBKSIP+4OXXm3taS70iViYmrYhWtKU0il6u
pJ008WATH/NNt80xQc7tji5HkzFamG1RKpX52ORZHu2G7OkWuiaZddKd+oqwEhCw
OkvHrtinyehZ3gsUweHkCazblCjZawcj724+OHen9eQSjGFkyVLjoT8sge7jag1n
Kz5rPQddyqPPNJa/6WNpwYoBrdRLZUuLRDp45YDreDquzg456lC4OHsOyjpIpBx4
dJDO9QOZ5jVTqsakzjlTpo6F2+AmN4YC+jQGqVjjzKefjASQM1cnyJyz1uJSDCMA
nFaewQ8OOp3AjQ6wM7Hg4YlvYY2bf9qi4Bnk+EFy09A4z+TbxsnZmvi/4mdhwzgC
4kDGrw/3B5jYg09U+ZnlywtLTbH3FZbtedPOkg3pJRL4ETA8iG5KDkHnMGpsmAuZ
cV4YGZouqEE3Wdg9Z6dia/peyZheuC335110Cy3w6vztJIs8HyRlemGI/hFYlroN
pnSdSJg9JATEzaKfnCzoZzzyCdFDQ0QfJYNywZlCsJamzYhCtSUf7c9crmVCrP6C
JJntFJvgZ882f04yBaznfllIS9xX/qSJ8jUZVRJmQEGGxSM8L/JQQ10FouZDcw6H
FP0Xy43dGk/9w/wX2+S5eEYL3XhTQ3ak5QRx9wgEGeqU50NDf0iCrVLUeRkcFjvm
/+jFcCkRhUGcZZEyEWRA2gycy8L22mpGLxzkAAk+t7GNuRaoZ8q1wq4r/dLi3HaO
pCOUaSq1423Hlw3UGGYvOg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HYJ0dAvSYBLkdQ0ep6k5WmwXHBwFiZ+rhljO78PkZFrEyGUU1tYWrvFfd8FzioAR
rnty1fGOkqmXU0lrO7CL+6Ct7ZviEiy3hv/7gBm0Cq/hmuT6O68ZJbfZ7+aACMzw
8kBt9GNNH2fF/WTkTMi5cr2vaD0ehGz1Nc5DqzPOYAtXqD/tyZJEpdHxX3XHlb+d
YFKwAcuGThEl0w3a5BmS/+UVpHGzvJbKDq7OgqBtWDorJUYaD+TYcY1ySDoFmZDb
a0p3Mm+71PFREpW3YJd9dF1LatXc57z7xNaDfYRqVwo+Z7cfmFX4oTgahZepLEeX
c66y1HpMGaOcidNh8p9Suw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7408 )
`pragma protect data_block
98v5F1rahP+/aaKlaDQkHT7wsx3osypXTChu173ITdxsYeFzZPRIGYXcF4nOfFFn
w06dlYpKkHP4BuDagMhPNXgp6k6CQpHcqjObRNjcxdBX5NFOgbDz+8lnjDsxk7B0
LGeDGZSL6mn/ymV/lquCACj9NmslOSnp3Tj8NPl1+EdRfsycfeDlNwzdkBrzyNf7
EvskFdLCQ/nYdCCA2qmGnbFIn3Btm1KCfekPh0/BOBQvhsrebyVkqfP6P3VtsJHq
NjgLvcg/VdvgrVmlv6FUDYdnHHLVjk5ZvBwizNsR5HZLM2L25GltT2WvQwW308HJ
013uoOlf1Baw81QzTFV/Ng/zqiDszK363KjgBt/p20QB1f7hr0hGescwSiwXQDE4
wx8sJV9SkzRNZ+ORwXJuxh7Re/qxIvEv+xGguYeiXUjHs/Fd9qmR+achQQmGe273
01TpgCPmE9C/CkMKU4h72ksWYYZnYC5TbiqZbEDyYC37750r62VROTs3ehS6/Hn1
4hy6g/GhBhrT8Ntkf/W8X3yR1ai6OYwa3O0swkekSbGawdklVfHO9wP4DUE+DqMX
Q9x14mpKrIqrz10Gm6l00UW3EBp7+rPAvqLDoF+k1VkdWjQZXbjdjYM5rhDBC79V
daeLQai/KOMSy6LPHN727g6yv9qe71pIKeyZXlpZZ0vWjIZxNt+dj5NPPn+6gbEt
L0rSNeVw0BhSjpAJqycVkz26aEzCQBsxjJxVk1k4A9hIFn5FDJU6KpocPZh0zI0L
Q1/QWOZ3CrX4kRwW2MRAFv1QmYhUYzD2ZVEffKHclG6xdm1Hejof3YvKkYpHU34v
nCKyfdgfrFT6Go1pIUmmQ1stGLo4jWwLZQOVX0qA443nK85oQSAdjub0G+okuHkb
roHwlXwScC6T2WOizg3uK0jehe77QjeT9I1UwYzu/vI6G/SMKnLfRMATo/XqHXW1
kVC4BW1XYFczk7odZgXs7/ugE214YzXQooY6eovyp7wJXDrQ60vGLIoj8BWsqsVK
n8sgEIm+wVCzUeTUEATpmZeembiahiNJfm3T19qUpY3eN3KwfSmhQ5owjfBoG9/B
t6/vCSHVmEEaeNOV0U3pg5uXOJ9xrDU48YXlm/jn7oxsyXCZWUICpdMaEAW6PGI5
gaPNRbx49RpL8TVSpD0ul2EAjKLJtB4HDZu3AKLiiqKtFIct8bJ6RECfVNq6E+jU
DPjXpryER5wYzbMoabbeZArK+WmcZvnwEmMkrI+Tu8qJSBAsXhVEFdMf/XioOhVH
a9n55cHttpo/SLUUBGtJ9/ymmhmZo+dwQMamE/zHCrg87H/mPUSJA9MHoq0OBpDV
vJwhQaHm8/3zcrtlzqjxqLI51GFMMiObrc4+70LkF17+LHLPPcLXK29qIX6ak0qW
D9goU+ApjO7i1WR/gX8nn1TvfMrIexXZY4i9edYisLyd+e2uJtmEe8Zg5NxL/kDz
nnusQNj1sFP6TMXVFmq2mgkUVC5eN+9Ad9CRoT29jwMZuj+o0v5P8zuWu5lZxBn4
OsEsUjlkoFrP5YXE2V2kiQv8z5PS/j3+26IWZx/cB1Du+9bg0/mDYVkajJfSt0YS
6aAVEXd0lFL32Unxz6dNPGtLIRBB7Js7uou+LIUmLtMcPB8RO8xLB0juhVYBmxAz
f9nE6BVYLk/dExPfB+PCmsFzDkZTdX7HYAb7Ugoa2m7CPVgfC1T0dzzhRskYN9QW
V+Lw65pZjVhJxw0alht1PJ/sh08/8qooVyHDB6iJobyJPaty1nP+qoOm0EQxjKd4
wKaL1qLyIFQ+6FJU/5Vka+MR4XeMcmuSI+9A/4XOue2bcBNklZCZV7zwH0QMZM1p
5eO1cl/SZdkaiwmUpDzot6gJEDyr7mwFuHOrAMiEg0lO6icKn4j3+BmP6xXhmugV
4uH4fc/N3og0GDKOA06wMzW2F4kfMeKmmEVL0mITqiXRcljqudUCC+ujk6ISB9D0
LJrsHcaVzRYC4w4kCKYuw4wDxOraUhmmOKopwRMDW6P1PV38gkHQ+nq/0DvvIOQB
ghrFu3afqrM/K6SZ+3wEhSCEx0qOWiLtOWf5604pBcmDeuzqTaK8c4S75iSrQ2e3
vCCimsSDFXLzCWAtfzFJ5NI4u+paGFQk0aAAQ0/PCrw4IfM/4+lt8/xSdeh/tAg8
+7ONQ5M4rPb1G3ThK2cVFsxsdfQjUFTfF4PNhJ/roO3iufz3FMj201DwuKojPgT9
Z7kIbMkZ8rCgX7SllDpZtjJmDrZYNWqab2CxERSQSvxE9PXHa2gTIBEvmYbey8vu
hnDzD3vLDnRN/FUbzYrYgW8cUvxeGe0oyBPQ1x4VbNuVBohNDfDmz1UzNJzsRDaS
+1Xhr6Hgd3Sv+RxzX113wmmpkOZ6WfoLofoS8Reprzeorgrgw1V7k1atWLDV9Rtl
gnaTawscdVmfx7Fgfuv8QylpvOBA1ew13ohKX1IlaRhGee6aqQgpJj2mxOqZ2kpN
RBy9JZN+oD6yVG1Z57II/9ureMLNrBGApkYyOM8Trsw8KeiRHgCBl9BPH71ym0WF
u+yO/fwo3Fm6M5l4TYhIpJWwhUMOBuBFs5sJZWw9nMZ9HwVVvHMkm0q0XjDWo6yX
H0s5ik+pA+LCFp2dtlYR6wbHd4a9wwKHSngN4J3J+d2jxUNL7QjM/eHBNtLVVHYV
e4KwAD9Crvb+3I5ic3GnolrCswph4f6RuKfSNih7Ts66nOFJycpfFEbfM6ld2jrp
YhZFMxRbeA1+UVyd8wm9ufxZVsMbOZjcFA1GUAolj5NtJaH9OkzKm2804rmG2347
oXVd5oPqMPffID5jKX6QvgpRuDUnEgC8LrRZnWOIQMnXQfoTO1cnvRNlmzHI1N1e
p1gNayFtG5AWhlYJZbpNYutGeRABb4i87A3rVHlJqqovpVico42zb+EzUtux3NbP
uHzu40KRFN6zkLbpzacMekkYJiOkR6LWtWQ8EOjRhLFGJUVFeQdtmV+om+Rl8Nut
Nrws3HK95Q59qPpzCJ7rJbsOrNPlwOgSCdfGPVDlDHWWeKh1LSjxL8UPUNIwYVIy
KJbU0/46mPfkdChWcrJeV16TBdOq+ZNsTKPH91GM/8fH+1+doD4829i8HaALLUuL
deUJ9gewfPR2zpH1e6Sq9VrylBhwVzxRIXypyHx8SzqHVzRYi6Q2HD75jBeGeixI
zK1xD05NS5gRSeOeIEKSZTk247dLF2BLnv/xwgyBCdwTAjIzDqwwah/ZcR/pxrGL
g2AnglBcFF6W0KlZLYKRGp2EVQhm8UkpNBG+MkBrWp1d76Z8K/TLeB73W9nyIZM+
wgfEFMMteiQKsS0UWQgSDlEPWnsM01ZNRkXZLsQoTKGdi+tANUfVUh39R3ZOU1t3
iFZKwQhIjOtiNtqWbnq2MBJw/oz2SMKePakaA9wJUt8FvYFqW7TpfzFrmWgzBlVR
SJykw/+kgzr6rYrqm5v398Uqd9Ps/RGHaePMNlHXNQYEWRNidctYa5W5v8vDZVya
NKG7V4NDEQEsFlQQx/CGg5GuIQZA9ErWqU+zpiZ9ovFnZ7nxW6MQ91HsF5QUq6T2
QQMRABPupkpTCVx/5eh2YGcRb4prfH3IV0tSZEX2sRthpAFupl7A1jI3NIixdKNk
puCXsAKU60Dhy4d5m7aefkktwE90+MqH8c3e+fJpuoAuPfDEJ3G5pIOAOsofIsFf
W7c0ZJnPJHI3K02TTVjyFpiF2A7zphG4WKUPckeacvFtG70LsT0vHLXhLXtk/irJ
S5/FAls+e+gQ7UtakLUJyLdseB/kT1eXdW6epgZr/rXZ+zzyFboQKSFb/J83Dq3o
KcbCa3qGdj5WMSc4+AjNSOmrXisY52Tt/Ra5LCxLWrb5qL25EciSyKjkUeNrwB4B
Vg5hq+Za2JHEkbkkpOK2OJrO0wx6R0r+86qrshSEy5XyXyqD2uWp1UNQtn0w7Lsp
xeyiSs9xGaM8+A0HyGf4Ex/KFbcSo1RXEaaNEFO9GP6U17dK3VsxukxojbInfXWy
N3FeKEtz7LNN3fCcFhv6KfabkDVILLz4epw3EnBQzc8mCL4jatryR4i7IuoqQQhY
M811rojql290VWpLNiKI8VOA7vR9UdQYFrNO7TxLt1XcJYX+XGrs9mwoZ4j1voL7
UufHZpgSVXuPRv7JlukR9F3iSumCkgaNIc/s7soHf2iz8IpdKcvA3EcDUqUjHglo
ERLoenMOsiq5AQGQdT8pVVQGhy61X2taIdpRW5CrF922jn6kKTp+aUYNCLrqxbOC
W4PRiPZ89VH98wsiokTMLi2lS7NoYAaAmKubjTbwv367dm9Lrgn0tzK5Gs//w28S
0qRgQCcBQgR7TVWy2vLYPr05UEgUJw4gV/kSejfa0opcNHNMfvF1lcBvF5e/O5rp
7sohk5qE1TjJxtBSTRD/jKp/Md8V7GKy67jvcQsXvHgGFv5t6N+ABz1u1cf7IlL/
fK6RyO7O2eB7XLQhy63lRoFBcHcpjOqIaLD9uMpbAx2Jkx40sOPLi9DasfUVTIBl
1nktYrBxHzilFi1OSt7cpxevfILJhDfsfoXvaBUcppshzACrFlr1fELx9UTgbqdO
marUZ9WqxUSQNYSAWI8hhlG/JrCqQrSCN1cFTJEqEH4QLOAdpJF9sswpRxPReZSG
r2BHwdb7I0gTMFDTIAhi3qwgTr1DqYpNXk0wCtM2SgF5ZWI0WAFLyV1irNpfR8AR
7XdjV9aVsuDPTh9v0LJQwhxKPI6+WAeTsXE+32KlxIeQCffiZtjfd5AvHVpIdH2x
iLqmCmtbEr8IrKyxu9FxlyUj3k+E1THaFX5GsolnH4KcOj4pVOQL2uyevetSBgac
0JM+r1zHEpKK+uFLlyyLeXvE69nmIRtbiCiCws3dx+P6KVrcv0E/MFUUjj50vB+3
WELLErPynyfMsi1v+QukTED2i/Rvi2Z9ySYPubXAsZO1OPMpHxohGaD+hoH1hT0o
DoP5L5YsTVFYgOdcGo/Bx35XN7gykRhF29L0k38NP9sREFtEPNoGqv9Y94IN+zPk
1aYOKQWwmbPRTMt5bcEKSQO4jso/2FAA5klZbYXIzJRrP5y8cemzOKZ0lMlwbnZj
TRHdYxSgRmOFlC7aSEK6thsAfGnUEu+9M97Xmw2EEPrzqZh5nctsWn9v2wTpnuME
Mjx8TTU4/ovM5lDA3V7NL4hNADfgHq8BCQFoShBylpUj1dTLiVRTUYp+SrFz8UlQ
xUi3ZV+U98nRyFAnylWiLlgOzlvvBQTzo4kgsdasiFpAADvfTMxsXQfaflO4UE5I
2t6Uwk54GeMur00cQHOLpwPxEM+DoP4mQRY52876NNe2160XpPpSr0x9PCpYqWDM
oiekAhZATqLCTPXoq7ye/nhej5AE1M0ZtZ0wPMQDT1il/WEEnNGj5vIz3z719Tn2
mLxDE+YJnhJn8uOWSAjh4j65bsB7QHi8RAeDq/pYvbbFzTLtO5JYl2DGTrGZ8OG6
F0Qaqki5ZyJHsgyz9vbeKXdtEnC9L7cM8j/132aoPCoEspkdLk9Foq5rJkZWW7MS
FR4rLLNEjS07zJ9oBu0VOORmrOwiMXzNtS1HXAJLPn+iSuN7OzK1+nQ2z43QpBed
CUMiCOUYPsfqVXPD3dIZmxGKmRGezNUZ47/KTrIlj0fdzJ+UW6oB0N6dSg/kXI1V
C1c8HqVfYMrybEP9m5eiNZ3DZ1FLegNfe6pk0timwrf30NCWZCsJ3LoSwGja8/u7
yTV6YU5J3Uov1YINdJYm608/Ev1arkwf5/f+M1PI4T3zqgFkFBG87Fdb1EDJ6K4q
cXzuyP6q3e1kXxjXabePrIcxDfyKjywN3bsPo6y7SRjpRzxl3A99023fkS9D7cN3
a/j2tcKUUR5EWorMp53DgSzeWTouNfptJTDzOv9CqMXnC00jmcBXnxsyBG3eqz13
mqlO05AfM7eXh+BYnm5r701h6TR2GbslxHyqywPj2zp0YOQvX63AHfQUJUAx6AKe
LHiC+aeQYUDp8QWVroAeWgZjnZ3+oJzJxLUAv/Cp0Sv/k1r5Zues7VxOvF8tcn/e
97thjbuWc/hjBNV7zBlr8S+gTNffx3e/r8mWq5ofoPUyced53X7QMHAynABh2viy
bUWk1mc6lj/F5vS6H1y1QFLZPPfog+E/+ypvJGVTNoWdtUDn0ZD9Hbl53ao0fuSy
G2qtbQPZQu+RLstCiGCiB6n7jeJOI4hbw2bAINbJGk7gsZH38+RwCuY6SBuaqsTx
/49lwp7rsHLGUZw2RhZeKSYXYf79svAb5x4wEhEhFoqhLtDHrAhy0/fdeZx8JgzM
CibGAh8bsomax/WpVvY9Xm8srjjqQJUGcxWc0iBWt+WKa2dMDkv/OYTR7196gtEQ
mSjQ3gz/D+cm//nqrHAQrent9wpdnsJcJu/wgDSZekqIzKJXE2jdhF9S6p8bNupY
TSDnkFRirhi3Hikd6hH4N0gomtiAzp8HeSgNlA8/YfU1gpk4me84exh1Kjo7CjIv
ekA6aIWQEIdEqFGAUQooh+wAzc89duIAylNlRR53wEJqeXBvxtKgzcfJ7pebe6N9
/eytfulqvwqY5BIASoovmUmfLFKwQUyCxhVTdCViZtxgox4KCY9rrX7Vpsqco2ca
fGhXEOwdLiP8T2pagIXU1neeX50NHwECg9Tlb4iQKbafUEkscBbUFYff+dUlqMMH
/Qo39Fk250LCDX56X3QLDLMl6RPspekYRlQ3VFIdNw+IMmwPBUPzrxabKcCtEYD9
BIL6endI0IdOUrgcrrQnuT6nmOKT8W7l1ayXRkrA3M++DjnvEGm84AxnIU+AYor7
ncf51UuVTYKxkCEbrpNF+gMh5mDRoM/hsPRvBfDN9cpAoapx1vCy9qSQGCKyOTKt
P7UXItiKpUyEcnDuDzFxr5Swrg18QHlazxkLBnd/A0VuHfK1/KObdueDxyG54to2
yykb3AMbboetmJ1vBb7DY/+P5f2Zpkb4EjWopYyBtwTjFO44GCXjrtEU5rpZ7R4Q
IUee1LVaKh04UukVfitUS3vyalpkcd7hWKabz/RCEInQnOacD2rzkHgqkjdU3qCN
D3t6XyNCmof4gw6uvauc6NiAGhTmtYS52idK2hPD3z9ZjmSgIM5Job7W25FMXIMu
QsX+PP6xLvEtEu7JtOGfHZjRad+xRRuqpYZsWyOsGCjqOGalnCfaigXvNRMFffHm
tjolay6pYgMunIQoWv5UYE9yp7nV2tEdOVlD2eAFh4NT5FlKXJcHoBNz4jl7bDQ9
1SB334hj7I0H16eDOAZouG0wKjRPPf54Rc0iCwjXunr9DZDg2GA8otlGxSjMzoLT
hjT3ri8ttHdZrpnC1vMxziq6lD3LRehB8aQtvsQsuFz1VTVTm6qZpup97cL50anh
OgmzAX5TioJdcvGFooL3/m703eEXb81nAFUd3l9oyFwzsNxuCJOR9A8BIwDz/Q3C
nDCFSx6N3uxC6fy8O4+L+5yXz8x0+94rDXXVcAgMrgrSAGmPPBxTSkxqhwacPg+7
6Hz18YEMpVLxlIYypS8F7TPjs9sQT3HIr4uDYMFdU9QaehEy7VLU3BTyJewno7/5
VZLwMfyzRkmsP7STNDvG6rFe5K0cu41DAdfMVibNVeDdOq1sCP7oEoEcSXDbttLZ
pM0zurOODod7QGX4t8Lu5JuTynXLudGISTJxr4rOFAQND33Ph0X+gIQzNGdW4b2a
zkMheyQdp7kE7f0tx6ij/V2oFk5ZO1se5HQDjsjnWKdJaPqS0hnhT3SfNj3tbaWf
DpugbWug2SqZIvXSUYu0wYuwB6pklrzVYJ4JtcO//27dyko7LczoNlA9qamtHWcQ
f8FnzG4lQkzaKNfpA/X6jYqyiNbQr0PeLwEgUn46yMTQb1O5Oj7pB0xW90BVqVK2
ceBid8UWOeOSPPa7sg2vjPRIPBizigwkVHoXXOSRubrq/pAcVkaEQPDZ4HEAVjc+
MKLuiKx3X852WlFdNTBt1Ht+gYd6APrw1gPzJ8HZ1L5jNoFAnjiI5hC3FcLqb5GH
j5D0hPqwJ11zIhGiXY2Z4eLCYRiF6Lbcpkr0JzWgBOJfUjN3/GpogI14+euK7Zkp
/kqNHKVOzhG6+30XmKRmGw7ZA1O03P9T+cM1zdEpzMNmaJQOb+UL+LQ5WmASQroY
ED8ubFbi4DykthIWuJzyU5XeE02rcQILTfpPbzqqQzzeNSNvaVz70WFm/UZ32kss
2ZXQyEZCkvwJWvqzix+o5I93GAP53/HAySKJFiBYCYO7acHgkLQVnOziuwWM+qf8
olle8H1NXjEXjb2LwdXqZ2TKS3jBmN2MwXhhyYY07U9hVnDd3aA15wlpMrM+CgxY
Aty1j8yft4ieyppPHmEhfMscZkxHrZNY7aDlk685Mlyup3MF0ONkyr/JVmV755MN
3dN0r+Q7D77M+7kQYt/abgWI2IrjuocRCWsZ8moSdzVNBHuNazyQCe85MX+pWeJi
kvwcjGBGAeUaKmDCbKzx9HPiPHef1Ep17PAYpL4NnVIRBwRPUE2T5XFPjnG0flGc
ZBBF6OZhfYCYtMaW/a0967iU1lygQeXlTadNqOrsBCWYE1Ud5V8hEGB1hGnOmYCy
3Mhmn0UWTyKh9lh8u7SnVfCSoUN2NRILlpYgcD2YQNXJ4kSO+U+A0umzAA6IYf7S
OAWutbplDhFLlO3w7YFiKv6AUR9v7dIXLOyTLoiYVmmvubnbsZGfmygu/P5vOg40
sM8r89xvm9POuFZG0dAASozQLxry7S5lVUsH+3xgnv1IPLfOFtej9+mqywZnMqQc
IehOYBLskJwLmSyFdZI7GoMXNYOKl1FFWraWW0RKENrlgpuwZl3MuUv4vQ82ASxh
jQ9BmavPSNWlaX3V+Dp5wKEWi/uuutEZgwW/J6rWFkKWmZeLAEPqYPEUNrOX3xp4
dkCDAeyJPT+kUeQb277YKkbZR0ION1HqdBET429XWxf33/c/T9IhYPzxnP2ZIZ9n
zOQcIZI7JHhAPFfrV1jTdVY1KqV5oew7U4QMWSaSIIrcRfFSi2kqMdWfScesXBtm
sFZvaIQgilJ2pzuEeVYmfh8ru4I90fuPXADeW0QgHHURW5NoOVF3+z2DCJq9sbVk
8l18h0B+S0BLFu/FVUNUQ/jiszokNd0t/401Vq69CzQUI6IaI8Er8pwBglGs+Msu
UnQ6p7AzVJznVwtPHy5hIdeiosJNEqXsmGEIgEEaZc3zeY5czugu5OAkI/6dLN3q
y7v6PioAGLN9H5Mw5/aMP/Hp+fSYjjoaZ1CndxDnp0EYoh5iP0QQqoVKktj163pp
AkwwnYn9a2yW7I/Wwdu7EbjweGIH6lLiVIDTkKCj3NWLOiYeFY7nkSi1bxis29HG
4IdxM5lw85qcxgqDotUklNdB4/mnB65b8aoUnCB7al+Rx19hxZGMr+ZGmhuVOFZB
ko6M+PDYPRWr9StwNX/sxzoy4XMsey33lxQhrz8CuqOEXkw3I4IRUD7e79UhDe3+
6QK89YwLOvVQT+4PPY1gLS58DIuuSEFXcBWR715Vu1YTXU6lUzOU5hz6VodI/DF6
qt43Hp+IheguLVDJjVafjfQ8MG3XudJrFCSQl2OANCjW7MLCJ0SmF83pZqtnQqpp
XVw2qjlpwq3ULfdXwveHDjzCooGUK+lA8Jhe5WSlzMaRP3kMoxesmM2/h8mg4Imw
1VwwpVTedQZqRGY1sTMx69FoI0tRJnlJqghU5+HmNCuwFqjQM3N0Qk/RtYmBug6U
sZnsLYZF7AWuJRuwXLUqP9QV6zXo3uJdEjCLvpeDV5niksFJYVykMfDbt05elK6z
i5UrJ3kjUKWRcEVPBqcJsA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EJx84DkxxqdJ2rzfIPUiFjStS/kS12V3/m2hIovbPCzYC6T8mO/LWE7jju1KD625
WJKTb34yFYi6Ji8AUTAiwfdkp0CtPrde+dTgiZxt6+FVYRmnD+A82fAyLyTiB0o/
0SWjn4IKv0fJYDGNWFkYbX1AiBQMuPHykCa06FVOR5+l5PpWRCcf8ZnNCzmAsMWI
ns8EqL0FUxgycKoLFsMIMSbJfKfyWdzbuZc3VACECmq80cTllyfnqqKWoBMadjXR
DGftAH4KYpNYTDyz1dcc93jTuAlEjki4n8X8OJKjt757hRwctvTzGi9mm79QJHOX
Pa4RC3QbZcrh5NS8jaXjGg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15952 )
`pragma protect data_block
WZr5FMTfptVpbV/WBITVvgJlL+Ae1W9WV2fQW76wGq9mnz1J1iXgItlPNEIajh5y
Tlv3YYL6oyzST5GhxkKMMOO8vucwwbPzrF6B+4bVG4mQj9kqJa8nur/gnDiRgJQG
Xnw1bVoxK4ybdgEkih+/OARu9VPJ+66KVn+XWy3lpAGkeubJq7ee5Hk3OKUzkbmL
5VlpCd7fUpAjIMUjJkCQ5CdG0L6i8vwyc8n3prSemTn8ptgunlhP4dOH/+YXjUOc
uOVG5mjlbPGnZd8lPg6Y2VFKBLHxA1UKbFzidwkIT/+0X2rp2tMOP1X8R7AT0Ybb
xab94f0KCQ2VQoEpsmuwYPF6t+nFxrncZZuuNYwDauen+HvPPSbOM/u1ovtFr8lh
Lta78PfDiqqOuagzaJQYUwOSZ9qx8OB85MYd0VfyXYPnw4hghbRtlLEdemNKSTky
GvY/V/NjNekSJWbVrbIvcKhrNZJCCmrCjG/2IiWDnE3KJl9dZM6GtCc+5ZUGe6wL
i5A/IvJf+iuhbmimmJe2JzyexSTE+OwrJij2uwwnRobBqSNWQc/qMJWywvMmYOKc
OVOCB5Je7ACnKtXubpg/UZ+4RNeMQhOk48E1AY2Gqk1vZwe+d8ylFWPiyBEO7QsJ
DUgIMGldbAFwOsK2OjyHBUm+8gOUHnuZsmM0s+DYEe7HWGet0zuf21pArFjYHvsN
b2kzcdBd4qYElJLQS2+MwlTOi3CyM3UXA/8+18JUCRe2piTyXqzDkFK26/49/5no
AiRybZXPykx3xoBeqY+CCNU00pr/F/rfv4c5Zrg9MqYc4RPAT6o3M++DU7q7/uB4
okELURNvBba5hyl54bWtUn6QqkyUnZdgb1NX/97Bln6PInE585VdnAkJ4RyqsRWm
2L+E6EyMOXEqNSXhvxpR+l2nIoya2EAnwv3Hyblo4Rq6gtXO7mWIxxOANMCtHGjd
/x1YH78rV6NIqcUpnN61vtePQb5+emFsPt049I/BmEUevorLQRRjBrjBL4SGVztt
/gnKctVQR+SPN48KjTYdDZSvlzUVM3+WUEfrDP9HUE5QBHnTnBjvlTG/OCPwGdgp
Z0E8A7V68b5pSfqLjrJZo488nv2/1Fnn1TWEtFhUiDBnLP+cqhoNf/2EBk4Ll5Fm
B/CbCd5wMefmEngAKSOpLazasrpNAwLg0oVjJN4pajaBrHIfpfMW/RC+/LaNehC4
NZ1obcaCN3i7j1d0w68K4CQ8whYTjHYWVwYDjPEMvZ/6xWvfBm7Kw+UzkrxTVQvh
rbJYN9+d5qLSJ1wPq9gYkCSRr3oYPs17Ntcbx8x0cBUuCLdNqBmIsPKWr4Ihf6/X
u5f0cytec67FNPcrdNnfi/SuvlhElUHgV0SSHnpPdJvd+IYgO86AYXtZYIeLLFpv
1Lggju2zy2Kh/Dygbmzth3N17W722URbXIkQV+OBL8yaF/MuuA3mN54FO641h8+g
kzHNGKpZmMfWS7j8Pc0h0oZe5F3wQAmo7DrAXwMUcTV+QsbOwaD5fc349OzWGOM7
Lb8inMIq20oUynisQOJIAd3/l19q3sYuTSiX4XBXl6urX2puWVR8Eqjd9kMq8xh/
P0BxjEnH13P+7hKL3HxaEz2ym0kx5x4HhPvWVLAlhrxl72Z5+Nf/0qtCPh/z9fik
EcL+Qnnyq6nyA3efcVh1s7y180lxkw4cS5d0vRhHsSpJfx20fgb2Olgmj69o6dE1
eh9vdB4/GqNacjmZ0CDn8zerbmB8zRuyA9z3fKf8xK6VfpVDhZsjNdbtlcU1jQKE
zZ5tTb/yyT+xcrs8vg1ciiNistHhb31Rt3ja+lPEqoX7GsQzLdzqVRxODCzraUs2
qf3Vq58ngmLOSu9Tztaf2TsaOrBFal4RWqSk9CdurmzjYu3u7M+7YPjgnbKPC+Pk
HADD2xKN2iCQXcvRY0st+Vst6Vzu7czmestmftx4cqAKwAI8wXMr8Pk0GQbQuO6q
GTaL2HQhEHn2BoMRmMGK0FbQLMO58RUh/x/8+cWcsvZNi0eg4r6fN0D3yLcHW9+t
II1Z5rh3w5GYSy5RpSW+7bW8JV6WooZpN73dRrf0GL01ly4gbe+xdSlgNMtReXjQ
UeRz/ogZkR2tiWa/YJecov9lxluq5x46jkRB6c+G8KQ0e9c2pPXAvWOoU/hcUUo+
lHFp+4HNL0bBBOdIgtcqdzXLuDGbTntE5P9mH6YacgEkMzxmn301Mo5CGQQm1yYR
zOayt+D5ixLgxnQ5Z61A3ir6urudFrSZgiBYeHjVS0agMCVtGYI5Wf7ALjmTQtoG
qzctUw2OhaoRV1Ig74LcZJvuRCb4hKDJMh75+IEKT+eTiZWEQsnJxeAYp4uAAvrt
wyKaYfNv6YvZLX8lOnDGP27xM0cIBpyLF7ecQMPQB4IivXuRKEg+/ipZeURysZii
HeGKxUwFtjBDnQL0OXZjMWcbS3k2+p9jlIV9+SIbNwI3PVhm6VXH8wADs0NjukZe
DEWbC9FAh6rwJTJFScLdnPzpkFV4ouBKMoSNBLor2bCoRkUjEw5wzf1VG4SNujNs
9srJuBKTUbU4QIbdqCn5D/ztvgds7P7VAQDjKZ5v6j12e6mhOHP8KQERX1pNxq6D
qrq76/OAYrCuNvwrg0Qg/RijVDHtzVNFZRSlQ/w/YuIIbqIeMucI0XAnx4PYJjYl
XNN2hbpOVsYCMtZ9ZMFyIPWRXHLtj5dLvNeaTJ4wJsYFpDZRLIJkiSzZAYDUquU9
974KAnyLExejyZjrJDj48tDOXi+BDAV3tAkOtWhBYNiiOfUFoGoXcfZO+wdW8785
ImNvvdugdY7mMsEGNcyceX2UhYdDQyFE8IPgWPQ7RM+H/U8UbvLCqyhgpQ/x8pwh
e6uJgknaZvh00IeBSCM0n04cjiyjFwXHfNl5QYzDySoMe7YGfBzqZ5PuPwYI7xmL
icsWe1DRnbnjNIyaULLfr4OqCOliPQxm0fGCunnwXE6RuUc6bRry2fPWpk9cUaCv
ax214deVAfxa7EZnUN4NTGToX4JldGdw+yV1I4gALRys8oc4jqxow4xp4Fv5cjLH
+kVBDuoJmcvi6hes2lON2Sc90FbUANrxYIV84w03iufJnN8X3xhVo7OsZW8vdS4y
mc+QY3rkEi5bDlreNOBEA+Ba4BQKQwyAtL29uMxOeukYTtOKAtjxg56lQTllaIsx
nX65vmn9UpnlI3sQpkXtrnIYEtc2FaW8sti+sxbwq4VBANLhzmBLEY9MAYvbwWjc
jnw5cyjqozOyiLzfSDJ1DSVHUdL/lvCz+wECNTMOEQADe3GagtabvRJeSOb6VweE
U8LOlGFarelHKu+hvrObanrcT9ErNJGmRRP7NKW7GGbS4R2/fI6rgh1EPit5C7Ml
N7BMr3j0yXKIYOrOn3nzVGOb9v+/8nA6VO5Smdop5BW30962Zdx5Env6VSXn6yUf
WSNbcIaaB4Zus4UiMDc6QJjCcqyqnpadf0k8i9BYlZzdF/OIb0A/kduFW9PTOC9X
j0in45oJU3dpTKVx5Bc4xRe+QALnqnoVWs9050eN1PbBk/3GZ44w9Q2phT3IEN/Q
z3pf5nk5HzUUFIF+S2kPoTPt8otAWVgh2S265FXW3/6JKS1ZsylauOwbzgN9IJTq
Q8rBeSSpad/VKlf+7AySTYmb4g3wrazbgqkDPBYcY9nTHS2dwW5k8CgyPJg16Owa
D1WyLMMWRYBXBOVx+AlSMghZpY9o2H8GOjdrk3MwXPsVOGyO5MRWWKOvKNK1QZ16
EcFiKojs/EauNelk1U5lZIyXqNXIELPLZbZMsAPdouGAi/k37gaOfuV6hX6t5ybI
4MxRufZkZFGz46maNo23wKP7c4WBPqjdqIwiR1jIVgcrCR2E8sqsBBEKTz2gkzYo
3yGpfBeu5rXshqIw4f+vzWxbF2OIjqBbpRUJ15cLGHsO08PUApmYBIr263BUPk6E
ZmplXa6q6FueSfJ233fRgbegpOem/hNQcO7OwaRYYGu4yaW97yp1c/ZFxheDZS0v
bAcVNyTqhSgQSmNTKYV0lK+tRVmgaowwviulMinkPHdR8I2Ml0NoSincF1xtTufg
z4hDSljHCLnvCXfrzEsd1KQ/1CeWKAEOchaJKgWicYygectFSy0pQONKVu+4qLzz
kTJSAQp0whTShXLD6cpzHC5RsGxcxFtqr+BU5KXAEOAYIoh9Zy/2xuiP0AeA8T3D
OwOiQW/yJKUNVmixGtdlxs/jRn1pkQASy6t/vKtgMHH6Z7qh9+J2DOd3nvYJyGh9
K6UdyzWFkEuP/yEkVgS79Alo3xJngEVmdgkBn6D7bjBwX1tWbG8iR1MO9nfHNiUe
N0E7bD9nkgv3G3XhHGM6YWi6hwagnFOEsP16s3rC5qjade88QSWydDNNHE6xVMXy
2JPn3hMItlU6nkMu55AkhKujiMulKLuuSN4hRR59bF4AuiWmcYrHc7FPncrskQTV
Tm1jK37s8eY4X+JfIyTPSvWGBmDrITCTloapdvYVB+W2/Ndb/+Rnf3mWRgmg1ln5
dbntruaogIgYpkJF9a9Os140L5+M5P+c2DFiRF8YuCyGnaO3D9uM0MYxnKoaEJqj
mBplfqb2pNB06yWc4/FdcJsi+r6Qo7IwJg11MEEoJgau/IYao0kcq0oKGdj4PfSR
k37cztytQUasFwnq4SxLIOHoZkenPqYNmJk4sSp8azEsxUGdDU+wOr6Gt3Yd0uZl
Mq4xtM3UyPVMGIV4rHD5S9wAGewvNA7dW5iDt8OqM2UZOBjffq/HrhlOYhqgDlcl
KDZ49Kz7vJvfq03ORlMTxhA0tZjYrG/0G1Xo6CbzGuVIcyNi6OpbqHs+0/dwrnta
OrWgWOTqUx6rZ1fXMvzhST9CTb0DQ+IUtqdMu7VS7ueLbrVramPRaBNkPsLfQnpJ
cVLWp4vmf/tTphYYy2OYMUJI6gFh2Ke/+Rv1hRMbrlRCUzIFnxJ9zSaXbcPQvcUo
bn4Paib41Hjd/leHeGTmJ/ALw2Og53/wJygMJn14o/KF1G168e0yR30zzdIgsC20
YHkbwXIKArZeC+a+9Nk3WcYnVLg8fgqmFQMbeobL9PlZSysMy5TNz5Jo+lkDM69j
YcrqDihv84ntN7waYVUDUaHjx8DjG13nmGhS2yXcECr/AtWr9JGU68HuVrQfPgDR
7eSApeW8Ffre4g23CnbnZGv6Qz/p0MW+dTz0mTwiL3iBoJ64b8QsRTm0PNHjVhig
gOVA9J83B2ubnN3barkczYyrxQrYVHcKnxNk9KZ0ZXtNHCryayofM+6HSrNg4Cuc
Yah+et5HNaVpwlzbG8asMU/AwwTiP4riRL66lvr4qW6tbk1ymslSaUu3Ic79iVWE
9SMUePbX7bNQg19wOg+l21sANb74t1sc3V9+TPZUJIu2yfdImhsWp8IX7Hu2U1zE
2SxGhQN3iH6TCKcVqqXuU62KDuJoaAlUpebgZjfI53iwNDuaJaulchm+geTgxknA
/GsoG3dh+VIK+9kICPbLnQ6rJGda9hd8hCAYXVy/P17vt0i4pC8w+/b57bsocdp+
QfMQl4K3nt+G4z2YZI82/+KiI+dB6oP+HZ/DmBInvbdr1y+NJfjH4XP6IdVVxFtG
5BE7rDDxFZGVnwn8mVbPwkeZbj+E25B0C13cxVmeezOMPyjcET1dFSlQiKAneuJg
sSx/qDYHKZxJ80EsCEqE3stFcPt8X/PNJVCq5Dxp6Zm8vx2sdWi89pNZzTK36F4E
ZTwXXveJ/LHT3guuLshB/0rEX9OOJai5MajAk1b2aUq3Q0n6hSIDc8+Mb+9nlgxZ
eN61dsZNm+f5dDM0yfTDD6bj9i5Z8wV7OmOli8OalJUnCS6xygRKlvb8TAiniljL
NWxmHMeb0tdA4rj1Nb6vRGj6GOivGBhO0kMFHEWk56fmJXPVJL00WFwGna7knD8l
KQeLnlh+x8kOmxmHwvOyXNrS4MkmdWYpPBa7K3ggs00qB+Z++9agsZO6wLROOWDP
4UZah1PYJyYGfvKvXDhGKqkUAoNs60e78t1NRiROCcGcOjDAjCn7AQtdcotEeXfb
mXbFQ8d8ITutbBs9CNTyyxggVJ7YuyC7uUU6JZo2bi03SF9vII4/qd2ZWdLOjADi
/hk3wn8ePiIkN9QvWLWrXeYOXBh8qFV+sDF1//McBNIeBuf6NGrsfXJcWRO8GBZy
DASgc4r6uxECrY4WpWI06d22GJ53pbd3UZrrSPbU8ETsYu9BJ28jmOs7SZQJQHSJ
eP/JJP/XISqaOBFxwXHnYjbiShLn7W3QfRcd6AXV+NZMv8pOgDRRnsC2gDnaTeHk
49Zy5qdBgYsL5UT8rPDbrDvUl9YHGBZKRxxet8ZGN/HzfBwtGbJVHc+VQTr1I1QL
fwC5lf4jk+Dsl5hxLkMN5QktD260yT5SPeqfTqA7HHKMcvgaC78IHQnDS0SS9Vzo
jx6UXClC/VL1cTVN9ECO3Ogae2YS8TdrcCyrY/S8nSP9qsikos7ydJo4qWFW0mso
YuFDgT5v/4qL2ijM20lhbYCHy3Xte00kvDBV0vNzUZIXqB6O6CEsbsCeHI+UFDfR
R/zMcqiSHf8Qt2yyNsFckgIlp1Q6No3xlN8uDtKcmEyH4q2vMH6rHSm7WGxUM65Y
kHHPo8+JDWubc+dwfX62e5EZptjfHNrZP/j6dgkFQqshda/NUIXWkPT7exS25QBN
iTZyPGCqzZFGCtc4HW/YztQjCmV1WLgmq9atveRKmnLjxAIDz+scEsaUVvMH83a7
pNCDLuFdrTMG5TNKoOBi/Zg3wPpZktXExwltQ45EIefWLS0W4ldYFb57QNxK/d03
TcshGfx0uQjU4EzdGoDnrrEvDtj2mgqzp02F/jNaUekIndfoKPgWoYD14G8cXrmP
o6CHHB2y5DY+YCjzs5vWZmW2hJEOq7uQNwTf7uxDEBf5BgP0rsUILER3OpHqUF0e
qgX2uiKzxU6Rt3knB+vqZzuDsmr9JPpVHICdssny0L9iJP/LadIL9ImVsIZ8SGP9
100mo02cI23uTE2aT0NrUkFYjBvt7S0D0zjrQzGyIvi0SC3xlNRklRyfMcxKsvhw
tmgKP++hKGbzWuLxO/eZr0sShgWtrtnwzLlSb0nrB3rEFaDN38OqmdPt5KaKMREI
H1iQ7YYfT7JqV5mvpR3Fyl26wQszW9BufiIMSUn8QDo1TyOnYh1tKcVVYxcfJYdc
+i/bNcKr0/9mzV5PmvG+hWLQpUI2IXBn2sh1cZ6tuo9vxQHGA2W0LVIBTnYbKnD7
blCpZYW1A1rBnB3Ne8hb/bLq65IGahc1BDAf1qFkjzBfomq9swwUR7RPTpscSKLG
kV48kIQ2Cp1WfIUysdUrNbZHtWDUCE9uL5s0lT7ehVTQ1pov7HM2eNLU0LV2y+lT
thd7RxQmYimO57dg1s8hbX1YzleOmT5/jELFsWnIB7rHG339NYSR4V7kZzSoxYGS
hnWW84zw9ounVjvEJmur9I2DtDp29bMjhlUYNEC7qPDfQc1GMtTOnOPD8D4WjZpw
8a4ixaiKAyVtccWwghCAVHqqQlm1GKW4Ww7E4ma7XA1qBq0L6Wja0lY6y/MLf7ay
iOvf4RdYD0zMUH4YjwpuL8pb2Z04+3CcaZ3GsdtCW33FGREpK9jfAyRXn6J6zblW
exNcF7ckgZrRBz9bCwslpZdfrV55bc0uKdMNPjQDadghBSn9btN0J1eLJab5yeTI
+ufPP8HV5HkI6/phTS2yjmLHNUeIoBcVVT20wPbsSp0Z+NtiXMV5Z2G4n11RiZLg
qMYr+7jET+32fxniBdsIBUeaQN/W2WkrizvhSI+zqd9feQJJibJ+PCCP6ZUQurp2
UdVa08zBbds7oeQwOdB1ku/2GjzsAYeTm2KYThqXG28a8DrJitq4DRYftNb6z1v2
klR2AZUHiol5fipy5tswuyQxPvz8ImxN1S/dZrFphiT4dK+jchzz3urbYA3gvDfy
ILCO9gYrGoeqZDXl3A0a7tymDwHi4IQ02DmPgMHr/rzZKvc0dZzzJ83527NdoiMs
JEWtRgChBriB7YrjFIxI9d4n8VKQVvR42OBBSgS49ibimPp7wTHKDS9ZPoIXdQip
Wcfj+XZuivo71oMs5/bxwSDp7JnZ6z7qmiXW3Q5ypTwG/CYjSLpb0kSXuVy3xTdB
nzQO594PejOcyFhVYZZKLOdsqIAHTT24a7ZfDoFwmPlJdiijA41kB1fKJIZJjAPe
p4d05OPhM0NyPUHGJGTFcUSpOlMkaqHXRd2g9+Ki2fJxeruEyqT014tvaZFmPdF6
jvj2tZIA1Ye6Z4lHTXHz4gdMKgazIS+Aym0Ulrq43Zk6HwQWXuVRdDcGLKE/x+ZX
NKqVP2qhpCBP5B8nIfdA/NAYAKrqZKS2lAkpxKndqEJEsIpjJNT/0rMiDj95q42b
P+/2bOMOAJQ3i8cXRsNVWrGSLrmnBILdO/D9xogYSYcUq+i9bbQmC/0V75Zc8I/Z
rx3lG7HMSRiDJyjeGJxvz3241YcHKXGljKWG4kQI9WetpNJaBRuLViJdjJ/AGYDr
rLEde4AO9G7W8NEo40SaL9sWkW/4pK1dIXB98Rge9GigWq+Pjkpo+5FJLwY4FWTZ
aMyTqxRz7ChTprVsWnPnFH3yiOTR7tBdgDu/LLnQN29gXHmaIAGxBYxsSpLjtAoJ
bf35ayWij5EOVJHXzWelKOIjXGWgKMG7iD4x3f95KLXwSbDOhays4i+6HVo7OnQT
0xM+K8FERaIEGrp4E07G5iimDICcVITFGtvguDYipWehxTe8wOqi8I/FvPXK6nL0
Ftneju+G8KUYZq21wWt9n6z1l6Kyt/bahD/NHtjwa8Z7i7hespRpeebIDOfgRLNM
ooOG3zTHI0GPJTf3bTfUUwohFFmwlzrxMWatYEoqccS5mut5tJLD62o1hXHFNulx
HdLHMyRbNxdLVmg3cHAYROuQm9izmId2Q+x0r8NKqLg8BNXqT0IgRlLJmN1FdLVw
W2P9hf/SYDVNZUftVKx7c5V86Wgv7zGyi/HFaqBi9VJoO4UGgNDeNWCWm/TI3v2Z
2PUCk8FH8jo2mTwqGEpPDY7PLdR+CI8bRq0mj9/TkTHT8/qxMKL6PAp0D8clB5Dx
2SmIb3XnUiRT3oB7KtUbBWT9wnVUQEBPmH18251ZH6Qg6PFq9vxcSJOjkCAtoRXI
L4/y9eL0oh2PKPIQABR111Z/XVKIHusm2DDZv+dqq9sIbBW2e6FGBDd1yb/nOlDg
RPGJy+9yBuU5+Z7ChTD1XZDXJgGrGv5iLb6Khu6Dr6IqWmvCNR4im8qJTewagy2/
sqLEkdOa3gdfn5Q1OELmfppTHIqKj8xRjbxo5jgqVyrBUTLhHcYJKj1gB9oMW38V
ggbCr3Cg51YW1WpbbQYJoeemRIDDrnH2xHst3BYDTGgDy+DxViH72eZsmTF5xpMF
FSqTMHAIB9jaxK60amfDiX9nJ4FCMCmo+yC2z+dC9Ceokmz/Pp86hTStu2YUztS8
0fDWTnyR9CDZf/ySq7ho29ScZUcZA+oqrUtib7SS6402/mPTIFTuG05qC+U8vh2u
NrH5AU4pXP6knyOJpLsYjokuAGNUgwi5lh9wbEMXbFvR4sK43oLWSu7FvCw7U3j/
ACQFKPLK914woLGDzyXnQADo+KNNhU7kdVT0AiX3PyhQ6TAovbNf0i12VzGPfy5G
icM8+jUnQ10nHcjTyjswcrc8kwrlagR0BwiDYlrlZWYWTyhZhnhucKCd0olUXvMu
pWW40/RBryqNZeaYh7GGpKp1vTmT9KKgn4RpHJphyfg78sXKS8RF14IIGRHeoV5a
gT5psWWeCF4jMmCcDTpUM5H1Q6j01D31pox0M2DRcyZATR1P0cxAq69v86iKUGXM
47Mnu7qxqL+Qr9e2FyA/oo+772u+mTvF3e1UparnuOX9DREEiXngoAGMCPEh6VZ7
eBh908WtM107VAjlNNcu0GEc4TheJ6INbH41Kdmvv2MZbteg2Ux7ah3j/4P11A6P
AfMa8xcdFFiXzo/Rs7wmKk1XIsTOU6i299HyMkCduVEfPkL62LHzMpet3gSrqQGI
fU098q7rYZXDlFIAzs6jD3fUP+PpgxBowOqJVusWSHNeo2W2PaxYtpLx3ox/VrZ/
2HIyyPW2JGQeqNS++CVXdYxREHyH6a/gzOyjioYlj57nkhEe3YVfbOw4DJdDgYL3
0H7HbXWm1VT4qS92OxInAAk2WKxMJWb2GUuaSHmV3LKsHOLztaaqKhdAjytXQ3TP
bRA8I1izvNFI5WmcH5R0wvF/2bkw9lGaRJ1hWaZ8cRqWEWFeTYE6UQW7My62GLOj
6zVEyyMv7ceJNXLn20WBjfGmFOl9tfNKE9D4V6dNUKtWd3YxUjUg3xbkfgybzke6
bo/sKyA3SnI41Eghei3n3ODPdkC+3uD2ppegguqwVRYpN+DBas4NA63CWBRl3Jvb
5JUO/Bj341iMkg3R7uHFIUoAOPuULfdnrDhqxcxue4naUyeHzbc9ubvSB58+4MW6
yoqQPLF7ahsgIHk8594zVbG44/oUjG8KtdULOV566kodnwJse+CFBkG1jmZPxhHl
FUXVZJskEG/Q0KgKew5fdpNBIZKWcn184NFuOY8Yies9Z+mKU8yS5L0k8yWgpgNs
BYRTgqBwjr5Qu494Ar43jPXQC2MFxvfeviBX1LDQjPh/r/usJ3aEqIJoN2iEYjeW
djvYuzVCUAJwkZUQsWuyluNgtFxXN0fH9E5En4O3CTnGyIzEUfNnIkbB2R8kl0DN
Uq0SN3RA1y6m/DDnJsPcqd8Khv0fS/Iyn9gCRm5YD4vfF+XNURJ/qwwN+YoHZO4G
tgWpqjH5pngsuDxi37j3h5lZr6vQbeMEI6QwOwI53lEgEh/+wnSEpx886tDONaC3
4dEeKGpxBfJHBflvOhBrQt5s0dv6FLDTN++OZ1ZeHb3KC384GBk6L/q8BGab5MVJ
krnSGidPKm71K1R9xJ2j20vuGbkNQVexrQmbkUz4S3i5t94egNdJHQD/m3eFjo4z
5XXWno3FlRmcNI4J6/ytRBvUOHQ/JhHPNL63LNQCUuJvgDKO4SZlf5fHF8Db+Ovk
5SKtU+kIHhE6T+gmvf6jLtokicUfbwXlUecuPxnWSnJ1rTAUJTXgfxHuATYpfqEc
Yv7G3Sh9hOOrF8tHt+m/27EnrR0Uqn2G+U4IaAw9KTMW0WH4PYU9wBQAHGyOIcJS
aVAM6ehdMvDj13Qf1d6uEriWikdqQurFPhdGusRB8qN+nOG3Oz8LvtYum8NiGlHd
JLtVUKg9G4BnoGqhMknbnOBSrGMVlcQfnAA6SlTxvIxv1ZFpQbnvm2pEAN4byxRd
EN8+Vd6negfzzTufZ80B4iEawquoSZgnfoUjyGmOD2ltYLWn6yvtDHysJErLY2gb
OuRcK0TgKwD+SEMjpd4Oy2eNqDXgbeAk6F8akLgu58Kc9L5R1yHeDvU17JqBQG22
TXTWLMvlasP5iP0kCVAg5TeHQSx6ssahJz3ZclufJodeYqDtPh+xB0WWjs2VmP4d
vwKNoomK5TTkLVzH21HSlOLNm4K+/AhV277piQZWu6wPLCaIVVeyxzYyRlJTvhsG
thy98Q2p2un/a0hOnfNQ2eH1pDggcajwjdYor08W9hMsbBPAS5+zdvP8RiyY59Pf
NsPYEX3Te/30/IayqWTyOR4ZsgNQN2oWgMwdMAHsuXpv8HjKi1XSHrYjhkWhl32z
Pex0ax0cPFzqIeIUiTrSHJNchecNNspb5Vilwlht8BKDYwExlZfyu1mePHO0nINu
ZSWE8ntQ8RxjWCbCTR8mkDnpT9VwUSnS+/+q5RSVX8exqmvjHnb8isr4PS0BPD+G
fatmQQTKJgyQM3Q5SHAck9qL9HMCRVikSsttexZiT0/Z/mYSYtAVyRcpSBTJjdJ8
UASRBfKsYSoWp9UO7tGY14FNIUfQmBFIpKkgpQDKSwyxJLYswjDBnG2Ey9wuQ+GG
DwhxNi1wKej9sNZdKYf3kq7iWyeDiU+Fv3OQard5W5y8UMKv+tQvAYKEV7DOc7p6
nAoSSE9rRD2s/nB63tQIQBu/MeY3YokLbbbjAyrStIBHoq6wLJSs9KaxS6EEj0SG
yCnO3L80+onUn1jJGI0hTVk1kW5FhreW8y2zbJ9YMV325KXtwgbQBlGmf1An7xAK
7SHYi8glmGoWS1HLOiJ83F9mtexOibN0y1mutQEQk4//AD2VNLmycPpBuqvRyXcu
A2K7ukL+KnxkunyJ+fgogxDTU8SkQkJvbp0y5eGQ5SeZA8OP6JXTz5ch2D1ucRiA
TAi+ygfYNWHD10QsZvuCQLM6DiiIesLDovQ1XCx4Eao1HSzguDDMW8wdvmf5wKyk
UQNeI7qg+EcZSpFAJbOnUFHZQTkhJBOy0eaWjctRbJJOe/fupw6A9BcudSTf4RkB
3avk6Db8HfCe2Qdu7ekCFWc+6KoZFs1d0qllIo54mWlS8I4t8fmEfYQfOIJGFjPh
hzS27RFLYYX/ilpEXcr1nvP0Mk5fB3y/x+acQVHOvoky0HXe1R9KUMUvNUigUsBt
+PEBbcHKcQxPisv5Jsp7TIgSBt7bsvedlxIwXBQ71E/b5PFvcz609R+1DbuKKgKc
9u3dMHrYCkpyQU+sVu9wxh5kwbV6z51UHtHK52d0Q7fFd1bUU4nIC+r+jQn4UhwO
YARLGoph5hFrnYwwip+mTeJt7pvqmzDjHDXj+KBpCUpL9iYrmT+wnWquwX6EktcR
2NRnoLL8muhhiydcxdmfTsV2qnlZ5w348AY7QayVw5SvlvOYzf8ijshudQBS5epL
hXFy/nFwAwKOYxBdX6ZedthNIt7cEl++1UVMVqri8MZeZ4aNlhcjNBfuYYj1l9xB
mEfrsehoGQGQhGBHEQikXavl4YzLVBu7LLZVu0dueqRAwde8Quyk/VJ1UJmlDp8w
V38iJBRkGokAkRTDh8ykA/2MRI6Z8eyx7iMXKXnHlXus33BvjKBrwAe6Cp9zwiY+
uX7T772/gSyeauHU5mX7stqvsq16WIbWdGE2naoc48it0G+RebNP82p9DtmdQJOP
EDCnsyjTt+zQe43KfD5/V6FNwmeNoR3CmEb3+cKQ7STD6scm9sQ0FTA6ejtNZhd7
cgYgCj0L9o5sXSpmmqJIDF3cB6/6tUcctHpVGtoRWzsshHQiYFTGr1bBLfxh6zhZ
OFMEh68cazSucvPtydF9AKut7tWCFEsDarDsyFzDubUB5j3kikGwV04FFAAj+nB3
GRj4JChBpngHwKENA9G4+l1L7ywRAxepIdLFm35uopUq8A7KkC6cPeSh8E4T31SA
25YnHqS+Tl07hnkt3qjprn/tlWWZgXK2MHfLk27ItCEPOIDfnRilqqXbyas2iY0Q
7w8h/bfvENKlFvJ14trIeW4+S0+ZxJ2I2OZL0zJYS7Oa+UY89foa1I2KAn20DsBP
OIqCvU/GUs0xVlVOqmLK4xoNRmckJNx3D9PbfwASprreJ9ry9wyirCktEGFqmByv
pSkC0eu/S8mIe1KOxk9vQirf0GEnFL9FF6x93dFDKPrMVfMCcDYapjnq7GYm5Ow/
G0XcQDcEOaPH9yXwIHRrZ3FqWk2dq505DTiibW3/+I8Gd/uDgBvhF/wUsSDgCx+W
MfbT36ckX7sL8xFfG7FOpONJfS9jxRA2oPYqfR0pLEmH7bKGJjw9D23Kedq3wpYW
O0sWcgtu38hEZX9BWEulP/6G2sSZF+zs2mojUUVALT+mIrEpZ393NafKo0/c+yrj
3jtC8SH5Gl/mOxf46auTLvDu42zTnyanGBJ0TGUy2R702vAwtwY5M4MV4hBtMXBl
eCxxTZoMW4OZ5QWgVizSp6+ua51jAnHka8FDcENXncp1SkdV4MY7oZu8YF02yfoJ
rYW1Pccud9hj6+2HUFe+ZrpIP+0d000s/3kYuX/vX2Q2HQm+b7YSZIpHSeGH5Dqt
kT5LkB34Av3tcd4zBkcQz+6eyLszjbfZhqltJdcMC3IN8zJNh8/diUp6cIdScaTT
h/+73L8sQaBqJfCp+1VDZCzfScvXm8AaDVF1m/ZRjZk39KcgPd7gCtAX9g2xHMQD
ItwPBiiA8AuwWF11aV3xJytM23yzlGMKXMef7iawm6H95RleMl0CNvgpl1F9hsM5
o+4/lZAc2nB6t/fgxdTeqaAU5j91rqTwFH+wFfYxLQe7yt0x7L7VdYBOzQ9tdc9t
YTtzQlpYLqXVoVw+deHwshwKp5Nqq9sB7aptAON/iRANuHFtXC1ffrv8bdIFWa3e
tsoSQXL2QQKs32hfu2VuPC/xs3f0kupFUyEdwUW9GKDL6RVmYDY5neSMwGwaYR18
QwR40+0TkjSAugJdRMQd0WdPejA3NtEduYHbP37fsWoPSRlmWOHT62SrmO0Uj2lM
FdJ/EwmWps69B8UPw2e3oyNDlIjd4D6/4gilwXk0U7DaRV8eonhSXYeKV7M+Dfxl
4xE6yrpiR5SdGhXwVtM3K07JKRf/5dnhq0Mvvyb66Fjt7LhvUFrtlDeUSVlIJTLZ
s0uVPl7ewGErjYIJcscx7KNvboqlefAYHo/C6NjvEVKZDAO+2o7XpkD2goqvbENj
sKgObFO8TUy1xkDfQ8SIciaAIJZFfipYjZNPjBwSdjIogHqqEAV38DF7JqHMsL/l
lJrmJK03dSTgmLcCM7lPh1nIT+yKmfMezoBa7H6kWKERs5jMtLURHoQp1sCOLM67
C+2FEy8WAHSbjiqBYqR7HaeIREkxK3HTNnD0aDqmToGlreFCjhR1uNCWN7azX+OU
Nk8MxiB20Ul+ZCNfzPBo4jPaOumkv84jbkj6DTiBGJq9TN9PO0opOMK1D1YoZF0D
FisIyOO1gYnuvC3T6E+8dJA7/tj/64wHjOAYNmtLNmWULck+d+GnC0D9IXpFGivb
w4uKdK2Vy4DQvoy+UdNfoqbwDZ5XSR0uR3PVr3GKlnTTjQnxyaVdAIQ++sGQM2D3
GZr3dONTMPo6kJtVhM/LuxxHkeUwD3ttlbrK8u3151WtU8G8WFHEJkQQN3NZz42J
aTILmqthXfBAnZEsDNij7XBVA1Suu86DcFYDVkXx8qrRVrpXygT6CxBs71Ksr8JH
CTkIdp6G9ehHQjYfY/sm959epaY5LacwvFjM8I/ACH0WmCia4O8PBLdGGk1rlh9H
RMwfS0BS0m/mZ5gdKRYz9egH31Cta7Ht3hsIwAJIfxb98bZ3zG4jAl1hcQL4fJTU
ECg7FZ7Hcxc1WmBAIjn1J27rdAXyMkCXqIQHRcox8ZD+CspiWzWEkcQRA37Ut80i
Yjf8hRgiNnb2CPMwUHoxYhn3RqncGEMM1XqwMKqT30ttnVn3ooHgfXqbyShEkL9S
4bvF4CfEz0rR+L4jjHPMhQ0u0P336quecKjgz2hIDrCp0kPRHO6vJ4iLKgAC58ZI
ET8fOZ0aeqea3NtTNJdzBc0/Cetp4zlC0VB4YyXP0pAs1vmblAAs/wk6ZvIXgBo4
jkqHIEfwEMjKLeY66rHYJRLSF4u/hVk/CB2bg48qHsCM3ZcruJMXH45gC+CDCEuj
K9+Gaq6dyrknwdTUjEZzymm5bYFiIb8VXXzQ/IX9Strf1x2WpTRDOhhghb+cNPg7
7JnHSzVC7cFrXvIDMAblmnzyeyNcy72v0bNgGXbNxhTIGdqcnMsvLOZPHN+/qQ4q
Y6yfoppuPkn8L8K9NWCXYn1pBQRQQ/BPsWRUMTjkF7vjhWrL/ksMXuCSOOVX7gqe
yT3+fbCznuA3tajmZD6aSM1XXPyaEiEtIybObY0gqt+fw8IlJxZf8KmnJl8NX2hO
tm73zIltGI+GFsvPS+Tk4Eb+INBAUe1XtmSzqUdSPmPeU4ByWE92DSRST7x3CKCx
AUcBECp2fDEm4OhuliB3W2LwEtWybZwOJekxnzMzfOzSx5lONafFIIPUs3elw65t
e1XrxIGUrncwiGkKJhp9fq20zvOoxr1jvaadTJKDR1zvbJmleUKNT/8Nsf9G8rDc
5dwB8FoOfGtWS5qFrZUjkSSNQIdv/qLn270dQtWVpzsJGin6Hk781LX1zYHPYdgJ
u8Y8yQwe82TIIAs/JMzF7W51+CQYEKSx2t9+tG0VUljhDrUyFfWLWr+spNQhWuNo
Te+Wvr3tMVKXDeWKgPOWwkjPx3AOTTrm2dGQapycfUJ//X3Gnt1Z0xsxaTDnuYRU
KDQt9b+20KZdUHKcrJ9tFLmTDMZGJpNkgvssptfbGlc5vqxM+STj3OgY0mx/7huG
sXlhTo/UfiZn4ZLcv5LrIyWzS318Fsj9LPRW9FpyZ6qtksU/ZyFCfkxr0ORTRRCE
YvwP6VRqcMZaCBsQCQ4j4jILN9ysQu2+SlKyf+nEr5aMJWAXdg0XMDCFnMHzyVzP
C8T/tXoLViY2s5gsszDC6Q6KjMMnoHpukyc9C+UC1iQFVp/6Dz0QOaOPFUV9Xrn3
WVPj7mJuJpFJhQPGMrXW3tIASA69X6cme/uUd4lX99SVH9JarhRv9tl/iKXAu3kS
5kjcX3efwefXH/uscAKMQECZycMV0GGfQW3R+It9GMpsHgdGmHpL/EE1mpCISkjz
EjVORvjyJJuTNvONWp5t2JkuLhxGySf+HQCpabeCiQamfy4wyLOfdCPSlrUbdkZ7
sW4ga4cn6AlTbNpVjlWTQa/XadPJx84ZuN2vMmC0BdGc2+Fh+ih51PHAqGZcri7D
S8KyHd1HOM9tKv+xiIu+k3Bd6GXg9TAXqwAw/3aP0IH1dxa2CY393afGGyOqMpy0
3o6jR8bJC9lqcSDfHRfUBOqAIwBn/IoLdjgxY8xLGAdHBD0rs5mu9QbMGhgZiTNI
xnFI19XLfCf2UCeOq0ntT5kBOS9gEKaZMQ2G0KFV1FMJX75m4IJN9KUcpCuitvzn
WDARx6+uPF6KmByOkCfmjJq1yHhIRBky2TpZACrVzdn/ze5GoS4CH5lzc1VBJZbw
aX+TzN0jeaXEmwMPr0m1TFo2v1XeYjDP3OoA11mPZb25NbUIlmKVNlj4oNrcjPf6
S9eymKq8wUxLHJO+JPPGNgtsIa93MaN/uDhcxmScILVa3rKVOaJaobQ+rmWrQn+i
3/Sr7ic80evQrWNE2o/EpqouZeyL51PgTZ19Y8IGMe8W+uTv/9W+3BSOza2YSJwW
0sLrKOUSNnPrR9ZLnOJxjziOY2d4Mne6BkisFGdSI4BbSQw13jdfYUseZC9b5RE4
sJZjU1GI7LBfXN5T1p0WI25Ueab00QB7Skw7owaV5PZZr58cakkd5AAmyIEOyb54
fYxWGIazjouGqzU5BRRqcAwlXxuEpc271+iFwYjm9fEZwS+DSKhS87s6PDpTbgeJ
z2Dr15Dvk/8NNosmryfaLDFGuvC9nnQ809gJOgSsiyqRxD0ZUOwhgHPnxcRayNwZ
WxIrpJqphMN5HIN64fOdL73ngZM/ZDz2D0FnNOZYstxZ8Rc23D+KpaMH37ssUaDK
9yesHkFs8+gVpULBr7unl7IV67iBOdSZX4+HwDJ7uYH2Ejxtiqj8gjAY7AgJuXzT
dbFa/rGxwg2PNvrxQ4mv9QI6V+ZJT5WWpMRqxO6yea6ToU8ZDfJMAt42zhPe5U1E
vv+uEJLLSV9g1yRGhoOC70jOgZpXyH3Xe41ochkQ1jJczySl0ZLv3KeObWIu+9gS
4PXfDmpLuplIx2ggoY694f0Yp7WAS8mAFAU5so7vOvAAzCF/OUuv6Tvi4RUqNsZZ
pBEoRvHo8+4yfvUbCVTMHlx7P9opR101Sa+vhqQRft7vpYVel4MNK73X7MxauaPE
ow1RV5Gtwgtwg8EGDJ0tchy20mL/5Rn6h3Hm7IB0qAKlOIc4W1BOA8CifEKqA2vF
QwFGPZ4XKYVMExkIhq52EEqrKllxASvH2Dh1Joqe+Gh34ieC62LELUtZjCklkpSR
ywqDd81Uud1KUMRtbciGMW2Ye4OU+NBlT288g/uz7I2/IKzhfAew7IgXENcYgGYN
AJhheOlRo9hN9WFT2P/xEnGRuzMRW2QXO45epbSnyWs6YUGPcEmmmvvPiZKLSlbR
oNEhvsu1Cbw7HJDHUg9dHqSg9oEbuTS/v3hplXBxfx30B0TGBHbyYNBCK7tC349a
aRGWDTzbHP+nwflwNaumuZBEXndeup7YxlqGPn2ZZw0BsBVhHz5H+ML0SbAKRG1a
m3sL20opTWpnjUastsJf41K3Bf9MJOp8KFElV5bPyux6YbrgktsbKUeaqTuhznwH
2Gd59u8veqyYL+kNp1qUgd/9BSi9caUx7kvwOVicjBzVDNaZ50qsqzDiGc0LESXi
AsJaY/DreQo2AIY67jdet1kLLLhgZp7mgR1Ci99aJ/xkT0XeDULaA8iQzFVfYxDu
+8hmdQIY8jjvD9nEClAOf7zcaVNHeCGdIyuTbk1edNIj8Xu4HAUTHdSmjHrSxd5y
K0/szOwAqx/LlwWpsE0VCsandiwvXv3CWepq8dezvZDRmukmLgauxsDUhOkSnfw6
t84p+DV1y2s8+6Q7WYoVUj4p6N3/lLXoRk0QVVXG+mpmmO3C8vN/adakMBeDmn1E
k0RY/yeUpBaD7ezAp42/qFPevKypBh4ZU5WtF1cYr2+ch2TyWlxcd4NpWVmUmlPo
wwrcmdLCSpXc+XjdxtGc22sFHoR+POp71J0ee2Xs3pSz/Ds4FaCIOCYQ//+1MFrF
YUpd7xPRp/Y7RP27xdLkbTzzBiS7FyqngbfnIMG3Gt7RAa00GA3EtXspkRk7Rm+X
AxVUBY8ZdomIZXqFspAoCmSWo+7LHnlBluSux9pj95HJ5UH6m3NE2oNhc15g5oHV
rkPsyvzHMMGVZ7LMtEM0JCXxaDo9RS4uY9U1J+SGYJqFLniWPj7QNPANVTlF+ryH
+G5aBX9KyOGlye45+X0DLKTgzYIpCoavWb/cfRph8JQUt81Zycakoo9JyNGWDPXU
fugdmo+Tc3Nuc5LeRHXk9nL1NjElE8MYWRxpuuynxE/FkzDOii+pnZfJBqRlRRaL
De7KQ69m11fhrkKo1XO0sQ2YENftWNHpJJSGPxLokzOvB994aYhexjZ16PRpUJTW
HI6VQJT/9uP6OtK4uD+v6HIuxclSZElVtpcMrXxA9a6ZGsc1lIvLMqk/GPNyP1uO
GxyNW7D9if03t9cg3KWW7qZMm3cyazd2566YfZ5P6NgCiiCVXm8pIuDD1rDy6x3f
8xUCJT2bJjyyVFua6bpwrJ5ZKugrBkGcANaENL/wZ9sgPhC4JT4snzBD5uVHuqgJ
i6IzgtLnK1d9rDKh8RmoGKio4BuIpZ1alIaXqvDRGL+ZxGBa9Whk0+KKdyYHde98
IgPQVAVMAcGpYWZSiwPDxF6emO6kYL8enDeag4QagbMgDSDDZd07wpo3eDsUmX0A
ujp45cAKqz6FjZVjm8IIpHzJFc0KXs51mgrMMLBKD6aP5xjHR6iGUvoKqDmWfIU0
es2tqA1cdgEa23Nzk8DJVm88kz/79spLMOOfvxAbCCQU+jaGWv3Lu83G+5W630p7
Vm2KmGXpUoYbA4iBdLMbhNjIyb7YW9L7AZRhcWtNm6/m5MUBNRznuLf7Yj6d7YDr
z0nxxbfwbkh+5Pk4/J7Hb+tMf2JP3evkXZjciutt/Cqxt88BnDajFpkhloFatUdN
71MhQ6l4wkVvQP3xN2Qz89dUmLnKFMKeKlKJ6pruZVfOz60/aAgKQeq6rrxrpcwv
CkgKW4ooFO1ShQ45ODayE42SB0jE55B82crd5h/7OTn5aMigt4Le8L8mwwhtZp57
HZA6b9YTJOnOWMWURpgcnO8jqRZf7akv5FKU8ZGHwSQ1VHw20rxma/qIJZx8Oana
XrQ8OYcZqUlO9KdCFWl243YdpoAYF6RR3zIa5KFQzEZBi9rwao/ekBF1IGrGbGqD
ZydG1wRpAabdW1lyB4x2Kn+lqnvc6kQF5R83DTLrqM3+8F/bRecHUPAd/1O6sFnV
xyY8tN5UOor4+j8nsOt/aWez9nCOUVhtEsehgzUzQeVHYVb8i1QpbtjsFN+/h5Wi
GQ+9N3xrV2cx3pR/J9P5OQ+xg7MFKEjNrV7mW4weghyDwx+mY8ViV+bzf+1VcOxo
Z/lENMjvIQ3KIAryrn07g/NbNhkO3/D3G2yWiWd8B52A4WRFkP8J4jgMGZjJwzka
8mq+0nRe38bdMegZxKHCz0XO+NA9Zhw0kDLS9aZlPRkLzJrkauvjxOe7GMHl/PWv
DWLA8KkhjXVQsD4XQLsO1gBxVND1Q88qNE25/6vWmfoaxFEgquD7NtkmxjOssg1p
qeyW7uSSK4wieL79udRuENJK0+J9jNmQ8rDaEl2p1nt0xWy/8J/tNaMhyl91ItFv
eftjTO0agVBai/oEKfCf8YtBe7uc6F5xcwGys8RJftLTjqOKG8WXSeCYZ26t20jh
VqV8RZSSSZmV8oHrG2J8IHG3LmSfokNlqT2hWoBuiYgGJVxPoScOAHdaS/BvN7Sy
Cgi/mwD8Nz2cJuBp+PMYmBLz5/kptZ0KCu6CHy6M6aHXhBbQ6gD53ncBpjCdYY+Y
+rv63xd1Lk5w65NDco4UvXNfw6uJ/Yi9UILfzUa6rfij027iJIstj2F8KPnYjOVV
TmlV7+QW+IaK74gxbjEwYZ9Sps9zFVWPY65hp9RLLajr+g7/2s8lWyAQcIMF/RjT
Y/BF09NXSDAxs5Oeq/9Ecg+6PNPXnzpA7dJalAFNKgTdSENrT+9iDR+/Y4qkmjDV
uc+uschizIkJ6M8a/GrPQa/5xjJNiGYqTUxoYV5nJvwOkK0o0oPhiHKF12xqLdC+
GDMIh9IZ6aXBW9HlvDtWjIGZNCzN/dRnMWYRK4HFWB/02L6wx3/JP3ZE9KmN+bZv
KULdyO265XyDDw5AkDbJYvNcZ9HZNLPAd34kLIp+8MJ6EHMMamaqdIlFt1E6MVnb
z0gxZOiZG38uN6GRGypbIOcwL4hO4newRLINNm4IErrGfZjNS03hCGUENMw0l3xj
Ou2dFEHerADt3/RF8Uq71gFyzJ4rvwRM4cSu69d9UkNVye3yK9Lem8trabvfHh1H
7wSdTqwP5fBQ7GRcRzXoowB84/1gKiRQMDYyuMleepOyeIwzXnf2DPVaZ6EUK7n1
TV3KL1B5N75zj88u48caEQ6QtwV+vBevoqBUBHK60ntBvLvu00ydOfaCJszGsC0B
5PEO/kq8JDUt9n/AqIYlDA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
arUTOjNYy6+Ph4uo2aHpN3OeokkIAh5JsqZUZ3FZH1kIGjT6/EIKmyRAmV+dx7j2
17a8uL0rJRKgptXj4MfOUL6WAGUKqkXuDv9QWdKYmvD7VtK8lpiZOrIZjKhEqk3u
KsA8+6lLqQ/4maTAYony70XglOgkM6paJf2mSA+N7dFRxDhkk5siSDhaP351XzoQ
2xTu/lUmJq95rJjd9cRH5zYUDk6bNFEzij49wJmM3ky68bjwWEqeZpMZD0aj7PTx
NZKPExVe+tEGpC4X461vSUocB4WEFLRY28HuWUWGmX8n8PFv5lhGvv+HNeynFr3k
qR15EQzv/UUKta2VmbcwDg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5616 )
`pragma protect data_block
OWetvGF/gI9wl1edsYxuAGkIYNEPyG6ilkCoD/2WdYhakTPhF4ElNAt1jfKtg5Ff
/U7B0g7jKfVgtxsYUGD3WFQ3dEhmQkHU/TWexX5fCBWVw3e+iliuITsNG6wRNnuL
Q102jZmEABsN6unWxSOC22p3UCkywDPVyrTvHkw21g06jc4MfY1RZtXdoHuBCjhM
YFTBNp8sBkLvkjiaxxWjSrlTYZlBse8cP7perJbeUSDLDchK/pD0oBvjcFOz/QCW
ZLZbKKB2GeqMswrZATxqTO0+8WfzzswfC+F4X5T4er+dlEYMAIUXRCElNnVhnRft
aaxcTwmhGkc9VMhmQeMcobSUJRxLZd44PvI/IxqZlyyT6R/Sh7LnDdy1UmbNtS3n
4A8wm2d/0PC4v7CVsU34NJQzyAt/Pd+VkOa1YK3WFQZan9ptUtS+qoxXpmR1R3UA
5n9MGeaVPLldcgMkD3m9hbSnn7JFD6K2CIcmDP2k9BzSnIxju7Gg+6MYMUuEepn9
CQ2Y9Vxs4COV537zVYrH14fgcwTG2CYqZJsB5kBIUBmCm37dyD6g1yCfjrnWrMmx
btkX3qzf1HWBD7BnqhFZ05dz0wKX5qVcSlDZMLxMrB1m9ODbIfFlj+fUuTZWr4Fc
4lELJkhs/T9agu0fifhXe6Cb8MnxXrX+uoOWeZEATOyr5Tli1sb+EcO+y7PPXa1Z
mnOIK/S9YLxPc86Nb5uLa41xIKc5rCPTeqJyj1y8xbZhWdSbpzLXbqZ4jIATvy0x
00jwXZqa8lK0ZjHwlM0Xz73YKWxLNh2GpBi38rGcthmbmbrrmPOOPxdfQKO9MBaG
Byi7oycffkoPJ+I4MnzI20QgcMnJnQ4e9rsZHI5HkuJtfpYeykI75pR6psYxfxrh
sK1w2Wgmd96Os6XF4hdPaf1+M2D7W5j4U0ktmobgg0OuMjOFkA6MtuFKCRzrSGLT
rD+cVTzaWP2vE60S1jyLRuzLp01gcNUPHPmtZauoN9rQCYU40YTqxtGxFw0eG17a
qh/5UqfAAj5NmSDS5Hfh+kEC17iI0r3Kq0oAxL+87IPFCO5qKxeCRUHZzt6k9VUu
Bi64shxdyAGMuQ15Cj9wUxiDhRF9FgbwRYzOs4NPcJKGebx9tzndO3mm/J2o27p6
2A/NcqKVTvP14dZg3stZR1kckTPHTwf2WQ/5gieFkxHM4JN3ftH6DQ0aMTyf9GmG
GdN/fu1aDShZIkA84KLNN1EuogyFFaf/fisl6NqFgJyNTLahEjQFuL3RUOQLAMM3
ktVoMYBvfukxjcpy0iK+m2CgUWfYM5tsAMaH3GOGZT+9SrmvkvT7bAAmm1GbW7R9
yHAu2AO/v+BvGKXC9raTbF7IVoq9EM9tn6vkNbjy2+q260mLVPcjT1olBxK7tCen
X//38pzuD1949zxpQ8vmzNeYAqofmvUvAb88GKfXQehIBUtxl6qdlITzaZB/1F1Y
zh0Lj7FQdBsE87ytqISDC9RC857GfkiZnB+Bf9SNKdebvAOQf7By7VD3+dN0CGsY
pKvXzcd5SQZ4fppVLBwT75AeSZNq9qHjw3oXgwokjz9Zno4HaNhhmtuAunc4GPtc
r57lRSct9gwBZpGQsNNV0Fq6DXm+s9oIsWea68wipldSzcGRb5i+ZofeKeRWYJRh
W6kK2hWEKapiGhsAgvdBfeJEy6nEsFunkc+rOZooy5vu9KfB/qFC6EziiBYZkBZg
FKe158rIxMuu1eSRptBgEvLFaxXoicOM7pw5hBmMoNxAj9K8AhCYWkSxQhxJtxuE
JRJXc5xUY7Jtl1u/wMwtnivRRpnNcLowxeSn/W+MpYaxIrlCwx1eF4CAEEPCDjb1
/jzGhSp/ldE+Cr91ryoX0EYytxCGjYqwopJWnGoFAPDjgzZyRSVOY45FYPdRT1M3
MDNh3PTK2UTuPuOUKdW+w2fjqaF4FEiTOUIVKp0Kgiv9UBvNr+a4lopyL0QXoxpU
EMD2d4vSuwHa4YkuI0BqwgD8jOgiDAWdHRzE1+g1mwFSZJ7yjOXlabiuMBcc4zNK
cXZUE1ASlXBROVKIeo5PWHXF/ZJsm4W6fo0GUOdiONopBcNDQ+C+qrHhUBYw/f5b
6Ps1Dy5k4sn8Ui77K71mt2amKmJCDTiMhy57NPACqXHV+BiRgGySDfpTeAQgAFqo
RP1YBXRFPdWUO0MHdeXN2CQLmctH9G6IonER5SG42dgia+eyJn+OoPedz5ycx7ar
todwA51ddJv6kvkY22/zQrA6zE8LQWomyrqcwzj3gK/NnvcCFWInWyfHkWfKlyX+
jZeNWbC5rYkRcouW9+ztYe8kVbQ/cbtMtM4VN/OG1HQeIC6i6Im0+A7j5WCCNhdO
hRvH8YDx4mUSpz0q9eQgOf5fdK/gyAzabnX/ay5qKWZZQo2WXLL9P0/bFqDkEWxY
PPx0SR0JNKDUudGZRPqB8w7mcXkAC2UI79lgHUgVo+6FeBWUAA6OBaSr4hVLnN8H
/6UlHAecqGTTAzc3BL7koerXBS4TRDNwLyLHj6tCQaokzkNvuUb1SvxKL7bncaiK
hrxLegCARFT9k0X/ez3ZNT4ZszHBERZ5Re6jm6KcpQAycZFZJ9ZtyUoQwgJRysO8
1Kvp+qDU8OxErIVV7nf0JEVjRYRh8TcKmBjpuQYM1PADU7VQrtxVxnXs4t93l1IH
0VOXgbwQVp1Q5rYyLY6f/HZwYYxyKHmGSozPK3zdlDT3nUax9e6Wkju12ePfMZmo
G9VZdAEVU/MOb4Q1LNPxpE4mcTPg24xnVNE7byrW83KPR5lUowxLKsQ4JfygNidH
cstwT+iZ6AWRViBpjpJ5HFELxfgl0cGIaZm9up1Cb+bYoyUn1EoE+Hxtp3Us/Rcv
POB65LxEX3YAbQVIOecdMevS92qMGxNjnfTCOEPlYdeWurc2Ib707g+Yn+tTCeME
xbXxSTy3GxvfgHcKZiSZOCWPjrz6N6PzAX814ATsliKqxW71Mr+VOp/808jEXiNC
MyNkIUK/QF49RxAeT5DVR57ebk7NaC93raWe0yhEOmXsSqleH0EAFhxm9t4G2TmZ
hwUGW+QyHMh6o2x9VTBO19Ow0+74tgEHK+jXTilwv9Euy/dslktb4s3bBYVS3Jh7
SZslkICDUDLHwWx+izry5CfqCyIaB2JLQNeRpIqElj5lPL9N6ZHMRi8RqM0fjiqd
tPsjvL1UGLVoFidefvoD0JItQ4l3W37fK7iOGtrVmat+/ywtp86r/9bpg6szAdxU
/Gpk/GaFKjkhkMYMbkUyXyYWv9n+RgIB+1iQNOPYyn3/P0Y2irvxPApJrrlQyCIx
K7up9FWmCjd7EQgHa//8/JKJB7sBZzddMYSC20Xm+4nXd6pnF4IT+I1uF4+33Wk1
NUAWqC/mo4c1bebgXzmujX6SIebCvlwMJHjckz+uhq8cvSFVclwDoRL2jA3lNm4t
jffc+FnuZoDel7iJ6DZJZy1Ti6dbX5POzH5vzfHoQzkktJZClY7Ip2cSVNBB2ni7
RMGdEycSkqqazwN6sI8nhVYbbAa9we3omtUEVLDWgkHesxOUOP0iVy5yIzuwd4AF
RDaNhmKhZFqZYAGBtQ0rpeRg3GvGmbuTCFvyw5VqGU9uTU2QJrsrEK9EMek1kBW/
fz3AGu0hNGK6wa6pkMSAVbbX3X66irTd1B8wyPMkMNU7RKrUdZICnREnxtgyuAZk
yC5ZzZ6fOcX+CW/cR4oY7yqnNs37io3Z9B7d7vmftEKxupAoeEDC6+pOP/DGJnP7
CJc3gKsawbcoY1TZLnnrTXSzlNP48oiZVppJEO3zPHxP7WYQJLf02CGnCXshBOE0
F/FdrmYhoJH2nAXjkTifKGbqnZSF21KFZ632udNTWQ1qjkLotjhe/+zMf8neYd8b
N+THRhn/VWHOzjJzmvu53Zb8cP8bbpI2wczE6IRwrDfLom9O9MrAdPW4aag6hT3L
416MwYqfbNUMKX0mbW/iqQdP4oEgfEW/Q86araYG8o1Oju1wOpzb+SSOX0/TZMFS
SO64/rGnld5LsrGEGJeYvq1C4tY9Wc2KuU3TiYO2HP1rbCxvW3vm2Y8NDIOENvEn
oe7mppnRZDbZC96AhsOoda79ObmihFVYHRdnuw9LHy1k5ON77UjXKltc6T1UshIz
SUZpES6UIC1eWRj2MWm6DqcnnaHPo5yTcUmMxllK9GtYUK1P2kFYLVoIyDmxL1dv
8SNvXz5KaD2OuR0I84V3FeXuvyIYaA75kmHon19PB0DhzzU+Kwiz6nCh8CpK5PVB
WCblQZ0TRJLA8QPPzhBYPxZ4fAG1QLEtnYrjxaqDSwcwsS+o7FEAjRU48nwFdFVz
of1T3QDV0Uq3RFmApdkbBhaGuRUCsB1JvYy0zIbFF88ycmpNFkB+e7Z1hcC3+wWK
CBarkxh9Ki/6Nf/MK0UE30QXksJs0s8lGoNQ/BUGteKxe8f2Eulu9Tl153BISl8p
Adratqn/cSsKOkLIWJYRDtYt48to9Kxr7ixR1rOGMrFaDNE7/C67WUB5tjDpBgfA
Smr6m1oXJJ7zzmhWCr/6b2W/JRvnADca0PQgweebGVSU0UVqC+0wzLNg0McvM+g9
EBWn3gZAzrU/dss3eBymjs3SJ5wW/P+Lwla0p11VxE9SrLVv3KZBFoZy8cogbh1p
DpWmlV3JHCrdvAYpnKThy5xty6mrx/04G/r6VkkhZ/E/A4xlh5DvmzjRAL91mrNm
cZAin/M6KM4GocExijxQpuOtN0TL3zladl7f/2onNAwN/la6QSeVcqpxts0r1jQ+
4vsrx+mx85u8NL3KzFXxB5NF4Q92VymhA2yoa1zImvwcNjF2mfPVIg58ldSMgzmL
4klt9AwUAmrPZ8xNZpyDR7wnuulznZTQ+zX67i+UVLCzTNZQxhzgsBEObbUcztbN
OtxHlQTKkmQQibNZlYT/xjdmDI25c6ofjf1A99ddapjQwciYgRnUjWClMfu+xE4Y
m30WtnW4peFjrQMdGFP6cBe6hnbwuUf+A1y7IE2lURkq3KqlCGNQOq0lMuOy6MjY
kuJfoIU5lAyHRRPHbAY7UgVjS1NVogmiA8qFWlUCOyPQ2yJQ3F2KZHJzYRa1TV9s
VfbsH9okqJtVUKH5Ic/Kwo/14F3Wv7JYjzQ0lvRqA6U3UiWRDvN9qLaYE7FV9aOA
3zaYsHEx1duUNIqPRBbo38W/0AO6el+LpUw/XTqoUFYbmVEp37Y0A5AInE51Emfn
7ICJhRsRVIkIg+UxBHvDIWEC4/ham1ku7yfwtIv3ebgr0G8tGgDOxANgQfJF8Llh
fxEUfBZ6KSPv9YwA7J2sAa0yyxtiJyldw3lLR7WQRKQBFV5dH6j0Zv6/1zoDLW+v
uI7zX9pthUjHtY/Dg/hFPSYIyzGQaKSZ7hG2Em0uF7MHGVBBtxCCzTdIUUEdo5OO
rUFwFRkuuLSwlNlDJ3XRwQN4QUySDY4Y2u6DDjHwMfvC9uA8y3+nIQh+LsJ9OeTS
Nzv2mSIbkNpAf8XtkzJqILqQ9VnnNAGa2sfQwU1BDoc86czIIYQ4hVXybvhmqu7m
tB7xLrgzEmOe4qtXmestCc909yatU++8BdvgaN8fdCZ31UYysIIqJHfZKKSa2hHk
0fnu7ACLn2RH2qj4YhOfPqixWzF99WLl23OwUTrvIHQCbH1wVzQjxeWJeWgzVXgl
Askvt7FsCxOkHV2WKJukv0/qyzrIVeCBTyITOiHP49j1MMHWF4YRV8t1yJhaiBo4
W5k6zEU/mz18U7uuX4fZeESZx2iFKN6PoXrqvaisLtZZVo/woJT+7bs2ZB0ofczP
PavCPOoBqUML4UWV81H4sk06+2k2oguJwZiG/cG/FIvcf85YY0TRHndkeDhAsjZ6
GKVuB0fpmp+DTlliQ3XT/VQY8c257O0Wr8b2s8RFXvpU3z9LGmhjTi08n6n9RmeY
jHn746HSoq4ZiFVvPfQBQOqZhNfKqrLoFnEoobXlgVJXUgeiJ8OaX6B8owjT4Bmu
Bz/78nA5DnoKFLBpCITMtcGUajRSAIW9O0Dh6Sn6bfV/t1jwDDq0oPs/XwBLcXPC
Gv2dXMbIlHbfbAWIIZNqKTm7IxA9DdSN5WA8Pa/i65z0egWpF2MU4qSwPGTB4VMj
WZBCRaFCvRDdDopQez1uXEdpdqpr+NImgoQbAS3USsUjnJ+OAPHUaHDovbrs5Osy
0A49sSN1azuNgrOBc6AsQ1AoRxDm9OcZyrUnhMel6c+vNpB6Gt7WVUy7b6AV33aj
FARb+e4YFat6hn85oA7TW+QgVroR9unK6Zl0Dul/9r8zHC/PvU1g86EDU+mk44T1
PBdcBzH2ooOClm2N8YfOLG/D6tSwlHfYMPIgu4b0QOUZYw8wJNNh2S+TKrSaXku5
qMgFdy54Jy5EZaHpDQyed7JDIeFXg6vJb4qKQvw+DgRD1hFAE+bjktDBB936AayO
s4b92uf8s/rPco7LrsKYPZTYv3Z3wy4EH4R4lFlXYXsHD8lm0R8ITvwqLy6U1RMb
V7b+dhvOBwCfrmJxsE5piXBXwuXSGkS38PQEm+5Wx9BgDHhMrdYXp8FL4JZ94Ije
4IIIKLJ/BlTYmc8rCGpUx4ceCzvkl2TZE8fJ6DGbX/zY9l0WriRm6j8uuhq9gB66
Qf3FMtJG44z+3p7LqZjOsjrMzCBMrjYZhKm4aPvD64oDr9uLZVi2beIKo+Pef5BD
nXVsvgIX0PA18FovWt3cbHtOO0MOz8kPzTvUUKwbRjqNm2Y7PLcIPTGTXcbZA3xw
/SZZC1ge15U2t40QWI4+L6HvVQWJMRg7X9ZSCzYFcaWC8tA0OypYeEMv6F5UatUJ
MeP7aLNIlJfIN/8d8rhgIJfiFtQ0nGy+0nqIfZ73xz1kAw/oXXJaosI0Oh5vAGA/
t5oZFtO7AdYStUnmv/yeuY0Fa6G98NUqogLngefKTrq5vR5HpyRqmPOG4WMJXXoK
/+xk8SwNITBWFCr9E3piSm4ZtDqBNRasLohCV+Fkxq0mtzRASnOmMYYOVbyJ1TfZ
V5Jfunh62qvFxONVUIOmXdgU/K+cNBWz6ZTJCFGElzLLaCux2jhdh1O4SZI76zSQ
IAeV0MapuzYq87v/yyx0GpCyRp06DXQAiPYPBJbTJx76rpxEma8lAcQrou7+gqV4
sUKdMkl7Ew2rDzVjhgz6kL2zlIjBONFlOUfDkOzq8o9RQyYO+oh+MhG3TX2XyLc7
tNopMR9yxnIFPVVbhASXTMEOMVKVv/sCt+thHqAWJROFb031E8wtkmwZxQkoaX1O
YS+VbHvLMSKuUbAEuwWcOZoIluurPU+ryY9kfFgx/w8KCMycftMSDUZe9xPXvyZG
81fK8UH9NRzu9XDrWa89HgvmmhMFlLOasr4FbZ2Oqe4SM1lKqmrZOmNE5MdMf0cm
UzDcTqXrqFO1TZl3qDppAKxfVz9/0DWJC5WfuNR2Mup9NRHmXRDyV84JMND0zrbq
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ld8B76YMNO6C39pGlz15j5sQyahEAJp+F9DoFlMDnXHONq25bcWLLvom6xQqtWCB
jS5r8r/vv9UVRDppzCJc1AY3Rqi/M42B+70ShXxsf9Pg+827W6ni+/b4qUwfPKAI
LQz/5Ao0IUPEAd+MNyvSH5amd+Vux5gUUkAo7WCLcakmvC3HzERW7eplY7S9BXJR
DribYBmYb3ch/RAvWK6WFUO82ZUc4g3RFPpbR8nTilJmSIzpzb170yfw/eTFXHgs
5buT2QNhU1P9K6+l/sSjmBWGi+EnkPp7k5I0DAkYc0yVuoFXq8BBT1WeZoc/Uow4
4sb7WBxzOt15kHHJqc/tbQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6160 )
`pragma protect data_block
gyLppNmoPbho5PpeedBQxjGCUD9+K0QcZ19OMgsjvU1T/ypSB/4wPIYVFZ6d9pKb
cUmQVFe/Pnt/le0jaxDgOQhRzUs4fX2gkFspDdMCcmmBppbvmww6bxGeINu5DH/x
8Z/VpRUEvo3z1Y8LU6/JG8y5LKY97OMBjUJe5M40xTLA0zPNwmiytkPg8D6SESQW
oKx4nn8q81u+mWftnfGATmDulyBTHm81uHDhEPKUqWLPL7vButnmSVq+0mvSomeu
ezgjv/R9T6hS9L3MDplzJfQjFJ0Vf0wDJY49IHXsAHm1H2gKNV9wxLTFqYo/Wg7+
8o/9d4ba4I31WJaBhmBnalljMT4fn8yYKJIdqDuLzOi9HG/ofdqFRHxVrcfkMjWH
iWCd0vDavYNZDwjHx0gjH6QHpQCi+bBFRv7588nTNG8byIVnQyQdEBUOBlzhcwIa
vfNS4wC222Yb57uRlsiVMdHWRIk40V1/EHFFc6vXy1ua9OMAWtnrLOoyvHyzAxBg
tXiG5sWk12toiEfgQBHXOaD7UNcBqghLoC+HFmKXqO7aJlXlwAihBQgTqmEajUSI
dUjm51ZED4rDaZ3s+zuA9yjz28U1y+eCzJbNTUS/0BbKKkQ905T+cab94tfxrvCC
wDNLSWRsoVYn3I1+c8byYVsbTlFJ2g3wuAzuJcnLBz4l9Sw5xoSXxPB1iYSR3yp8
RhbwdaRrPYOR00Bt/d79iOjHf7AfdUInJFtXs0H8sIoWP5wBkWZFQodzdEzurPPV
AAozutXr1nUI2WsG6vBnGV9lMwwR7a72QlfM+0VmE0JSWoUq/bAdfwJhLCaZ5R+v
am0rzJR72Pw2a6JPmoYzqaofEiEfWY/3pOSUKbgBybmKfeeLM12vYlz+5AIEPvb3
/AXjALRZKa1igfB7zO2ea0jJwiXz0Yt/FlB7MjkNdhkg5GGWC3+r4un3onIrUIjW
q/d4pk7S8TSj1S/H85uUc/JwZEMaIFsqcZcVtmHoPSD/ONqXm+4E2mLbLgNX4IGD
MT5hV28kcCtrTcV5mqeYmP3EVE8NAPAb7BNfBv76YdKtkbTGJY+B7Ewsx31XDmyv
+zLrheThNaL7vqGCO3E899v+3mTYB/3xHFYC7/gQli8RY4XwK3/mvklyNKn5tTkp
2CqPkuk+/9lmjSUix9qMOnE56Pv8Lx8Tlf+FFBBUEzs/kPSA0tLpTyMNgoHRmUSp
MIJXuTozx94XR4F5RgmzPX/uShxS3yVrWK4tyyFe8IHd6ybadStHYvbIZ1nPAz3d
xC1J1uMJrCl2J4GDs5wJAWRgU0WeUup6ZnI1Jx2uWMylLUi3DTbghm1qng+If9Ji
W3cSK3FJrISZG9+BKiyMr6kkbMFf1WhWjpLzliGR8YjxMT0LJYD82hrwztSVWHTn
zYo1kGaj9PQO9bBhp/eBpFvoY/MtSZxVM7sVWmsFQKdy78P9vWt+uf1sIrhMhc5D
1EafTY6bTnCauOPlgqHBXYUQYR5/WodGiTCmYuFmcGu75oSA2EzYX/1btpEbSido
yzs2xY7giNPMnyv8BhRV16Bhx5YZ1HTrjk/T3Nk6eGOYYELNqsDFFE0r1Zc0WJ4E
OduLuVBpY7j5EZ0FMJwyILrPgDpAwGGuyLMAm4qEC9B/L84i3wexI7obb5SMBjKJ
l5OtxrOncTbSGL71YhUi2JaNKoRKvIQXRxAqF3oGhrRMj0v0pug5Z4DQJ49T05xt
ZR7mC2KCTS5Y34rXYliq04LDZsuoLnwlxiW4H/zQriQjuGnU4unyZUJoIpIunLvm
KfwgScx/GF4sIjgiJdivCjiv2WZYshvm1N70wdMUHIGc18KbNr8WYO2t5tC9tLMK
edGpp9XzWky/pIFMnAN//zbE4wh1fvGVJEPD+JO5DBDvjX3n3lXSVed85Zu6PfER
0jaAxTHq2mjwlqYgX51JaeQ9OA9Yzgy52zNMfdClSJCeyxhvQFY4hFIWRD9gI5aN
ukGPbIfrCHmNvK6F32Fu6QdveCQK2tz2utXv25408b0PPJum1+XXFqN26mVMHZa7
V/P+xFnH1XkBF624Ionj/0vnLOD4bRLJak1DqKM+Gn1nByn/VrVTWG1j+nbVqy59
X8U5c1OnjpYOuErqu098XmG/1AIcYCEkasfHOHnPjpeyga+e6+3MRMmJ4N7oU4DN
DsK5hxlaUm+lpmicBXYQ2gRFzTlUEXn2vEWBcZsFLlzO6Uj5QZF2WwJNrBRnmhss
pSS9ljZprfg0w3NY1D3RL+h07ukeYjw3Fruswpf3naVnZaLRF2JJkZ8W+oMGPH9h
pF0KLDZk6tfsE99shiRsku/yFcqoU7KN85Jc1awFBtRU3+PfCkJekJzp/7ookG9T
J3na7zPbY+CsJgFKIDA6tBm3g2TC+SngDadfJw6Yj1pajFmrGwfyQGr7d8N/7E6D
MDDsxTN8ZLr+ZZMcIHcBl88UXcuRZGROveF8bJ04eZMGyxYZTAH8aYxTLpI0lV5t
1xjcmBbcQePZBaSM0e/uAQZuC9IbhLKBGH91STXrByS8h5sHTyl6QWkfDeWUlHkE
XdYztZwu6uy3Z2y7AhCI2FjYKQ2oA4H964aog095AWGbY4uqxjFZ8a5T74drdAuS
XZLf5a7UlzmKr9BR4AGgBDBBEBo3fGXuqotdWsCajDZXDZ7O3gKD2AAHEbN68m1K
Yi8506rXjrCu67lj5JWte53/BdagJAlTCw939qPVnWnJcj4Po4eKQP7hOKfJJ+zB
hViZlY55m/XtL4Vy6V6LMqx1YhBYk73GWKp3C6DIs8mMXNvP+r3COgvVrnSxzZBu
Naf+gH+hGRFewmzIDhGQfG76onWkA2Y4H7DiH7tYDSLnovHSOsT9QQF5z1OQumQe
JqKlI87BogJ3pz6HRk1M3DSaHKFUmj8iIkyG9kDACGhRaj8rKnHdevD06Vdi32X1
EdUX3JBQeatEcnrT4GJAtotLh2czV6wreEQDLxv1JHdZXCp90Tsj3CUMonWeZutD
zCvp1y0Qti8VCaykfQvhUNkS821tzx3HfJmDswnzoK/1qD4jUGdOp2+TZiH8fNzA
i+HtTelHJwCYQG04DBxsEGgNJBdkxKbFhOurIV8IU00bfW2exwOeHmhPhj3FyjN+
39HWo+WV3gs+P5FSl4DVJmVnu5SXRW31KvJEsYXoEcUufVBqRsHGAmswPlWofZJB
jhNg0TDp1c6bXT/HLDXud4WpoiiPX5Kxd3u5hholqhsbjWE2HCxHZ3HhJbi7Y2Q2
D7emMoWMKdtgRMpwuPppe6k5Lgq4g5LttHvCYwjVOj6/mEmY1wPsztQQnfB/osCi
7COWeQeQ2++Aa0sHUi3SXWxI63h17Z99KEqNLsfug9TywpB5F26eu5KUlbVl94s1
6xx4QUZiq0J9JJb4eOZAbMSsc1R3SmfNHY3DCH/crzykjiXYfrRUyCqJls9fLze8
5lZrSNTqYi3tl339qYLyKhawvhA7aNdALrCrhQtEr+TpJDKjED8NHEsBt6Pih8EE
rZymLiTGaeb5kDTZHnFeRCPyL1RHTYjO9xfKkR3XVrVZ8vuzPsdPS1cvOQpXTX+Q
vgrEg8OVhfgI3Ye8cfymoUX6iNw/VCbdCz6ksAnkb8Dl5IsE5sUtWO7Oa7sHHzax
UhiKtZ9ixd83M/bl+7UeE4Zp8ha9ieqQzTv1lZBQML+AoPD9wE/9IMNgxTG2Dpnv
pWUSXWIzsAvy5G79aSLaPmu6VI3NYQ1eCPZyuIV9MqQ156zGXiEk4u9jMK3sNrZN
mNdLvHTEvzA0PZywYgOnwyIUKfO91TW6N9xrFB57SZcK+9ERbrpqex5Ypmt5FU51
lcM+wDhdj4PK5Sq+03KIJLYY0h122MVw3U2AR5jjkSnz2fRzmfCbl8jAyIY5Q2nu
cFGWyJKwXekwOkYoIhkpAfuJJBfXSdQnN5MI/OpQSWgiuy8dO4h7yMVj1LpO4OFT
H4C1KdSTjNsYo8gRMe2nO/V80tNyQG54SH4pKdGQEIJANPevOl90qKYchyPpo88v
BT6xPSMR4kkC4tqyBO7Y6YnkVwO5spGpkDdvS9Ex5qcCE47+ArvXi/6AWdaBfy0Z
EvsnPZLIArSJt8pJvSi4B71E4ItsT+TjRttWGrX6HnAJ+3CJy3AyqY/i3emBDLDx
oyq9+C+jfgCj7hGIvP+jj6och8626EKnGC5eU9rJ+TErREhI/ldcb7JiQNxcQz1C
ydH68goanVDW3Qy0LIaA0UoQhzWlem5N3e27eeP5RmiMoIrkKEdq069uv9u4wXdu
in2xPfEN+W469ge/tCDEKN3i6qmTecI7SLtHPZBQK6DRmewDyw/P1ko6Qv8gkaUz
0othf4RgQloRNALCswlV7AF7ksDu2wjPxaxqbFs27LKENwoyKLelJLU4iC1lCFxi
Dh3jq0oyrhz9ZsmNMczY1Hh8bbCHmimm+fcTr/kv458QpmAYc7dAP0VWla4QLJhe
9JhliG7cvXknIK1bWfeitIsxmyGfwThAJw3nRc9FwVI1narq0Q9iVWjEZl2YcXR1
Rj/Kv81ujrb+2aDTVbIBP/oPv3ZXdxCTngv9MPPjN4X5PnIbmRXBhlxEsQPl9c4I
XywXhhL5+qFSfCEQCT99lj4Mg6B3u/Szt561G2zcZAuiCEuCLtQsdqhlM4FQPbCX
d9K/0bzrVuWydu4fNJhLJHEDbjIUq9vlHSCKURobdRI7w5txflUfcdI73qFpdV9X
DBhqBEhbr4NCUUxY2cWQEmvTuuqT64umk6QzMqK5OCqKd/BYEnMtiNpotUY3DgQL
Bm62Lwdu6oENYUM3ic4r1ilNjuCowi/TGE1K30Er1o4OF15fUZloCFtNZ3yJzZYd
NZDroYRf6Mnjj3axZu0iw5ZyJTnLQKOOepYOvuGS5tLSFE1tXQxlHMGkiFf+FDPU
CHOQJElOEAFLimG89efRMdwX9m6qqldTmh+NVUOBUWnIQj2DZN0uCh7CgwzVwOQ6
sVe6UBKwUooiRnw4LoLLxo7sbiPXx21xYxjvDwa4pzAPQUO1lHwjCCEokAKeBNoy
3R80Ertp5NYq6kbUSSVtzh3gHU93JqwmXFkP1EKYoslpq1PFMBKR6kH1yxv4Bk/c
gNwyMU06s7xr5Bxm+fuinTCFpUDjYFSqUXF8qYb6bizPjaUzXpWBgdr/R/TPC55S
Qznbk3famkLn7S1BYKqI55lZI9YS6ZtaMrv2giDHssCBwaACquob1yjShEhQHHj5
yRPCryKsjQWIIZJHLdXjuo4JMKCU599n3bEspNOAjfCkqBk9/sVPWZTvaGoSk0jI
/0CGuG+wRUWqs3s69LaMXebY8rYOGuF/n6eHkhYqigixm4OcwSpS565F+NF+3gwG
IsxR+ZGyGXZV8tEfUCnibZCqKNtvQVJG2Z30DelhoR20TmUXzFheGmyl0U5YTJ0q
juB9N2wHLv5S7imuWnm0dkdRiZKwGISlmWWNFmZHEXLyRWfZyqCzc3ZKgz6E48mP
Hdjx7PHsH6lGQ91WWKZKCiDlxE+XsaanBlIsKg5U30sfs+TNwb8KC6QOScRGsTSr
MG+Dn4+GAVnSBWXKjBJTRZfLki2MtoUGyYT/f7pQ0fnZ8zn+G6twml7Yr5G6JaQC
gtnka4l4ehV/M2eb9dDcI3W/xWwPJgr2dBLy0Zhjp37JhRKy+WnGCjSoQhqPXpU3
CMaaxNbsRyRafnqc7TTlc07/UZTvr6IRHGXa9nnkm8T3UZvOiR8X++6iyMz9ZfsQ
RpCRujk4rxfytrcFF497szkuI77eTa84Iyt3Bd8h+M1XrWmzyMi2Hv8lhFzhtE+Y
lFzcHXii8XNBnsoVw6HVGq8Slsnj2CNPqZJamBhylQl32P29J8uPLJiZD4cowbKn
da8ePDJaAVDwRk54VbpafElpxxYS7hhWodM/6woXI0tY81nB3B9uD2bwRYVWubnK
11YDAbYW1VMcO0zpX67OnT3wblApCY9UBN0PJGzir7Qp6tqlg7xjn34RpzUKz4Ej
wwPSOMNYHWBdn9KD9y6ssDyD9mnfxF4w40JYkxzVqXx0FTH+jCVInnNKMPkXUbrr
rb/5mHv7ZnWWRG7kZvMNJFljv7/tcQVAAtJs/2tryBgfgSJq7mbUtFoB2/1aCAW0
NQjH+or8UGdyQHUSw7YthMhmXzhfrInb9XI2zZfokCsGfbQ+pib/Kx0qpDBuorfk
GoZg9p8FcfnksA0I698CVTa3KroSFtJRZaRNeAzOMkXf1fQsGKtY/g4E8hYDCDAY
OITfDAwIehMH3UTDJOb9jiCME9iZLFx3aFd+EIj64liu6KFXyIBUt0irZU9CdD7S
kUyfLuMyvsITbpRNsIwDCYmjP2os+bQsIRhVpjkj+74qsQlcSTRtXiClN8rxurq+
ttbhbpga3wkXehSsUC8hH0qE1qOKbABcEyCRV7t1WsdWdYpyG/t8CtvPT7Edo7d+
04msyrW47J/9oL0XL1AZeHW+w1UhlgS5iGOuhehU6YS8Mnl3E1iXjCaRdQlxzH3P
Kf752n8BYbCyhsS3yPUSHDEFIXz8GRyVAFVezaVSLlIg9H1NUOVO2VcWLDrLw+ZR
7tKZELQv4ol/GKQq4k8+loZ2HN3DgkVhuLxv1j6GPiy4+V666TJvyLgarmrlMqqq
VWRDk7M+TfbapBP3h9aqYdathkLX0Hp2Eaq9LLw6lxNBDUZMsHmyl9A6QVOoM4RR
pETtVY3vkWkhZaBbzujvJbjFGA1gw7ZxTdfEvERFoUy18IW7n4A4t7QnO75AvYH5
4RDhleXdCC8SnXXqO62pxAAAiFMcDDPcAHT2P8QQdIg+ZZAa41Cl/cX3YF0pxU4t
/JmNxsRc3h/SLxL38dBflY4J+jbLKJ5K9OtjCH3HGMfPjk9+FOxoScwCEVAPOy3u
I40KR3Zgzrr2BbALOHpOhzLWmB//4NF4EtXoXiV5DZf63mdXyTIjd11yBhxh99Jj
xn+GGlo+F42nDoQt64fVSrSOnNveizi/FCTckEDmvqpXGhuss/kqoQ2roAqEFK9v
FzLE8cZEY+1E+l7yeXkkDU1CvC9sKA/+oHnfNi5WXipmHls6449wgbCDFTlk+W/v
OEDnqCK1TWeQHXTWI/y+9P0pgp3ohCcyP5DLzUHJlJWv84RvO8S0+gPOVexoypmr
CSDzd5m3zsQ87O4D6OtegWxdIriPdVZ/AnC3ylPArVuw81ij3oEP4F0wT69+PJqb
z+hExckkAQxGrQknPEycwO25lRnvoMyJ+L9MIq3WM4MFaKlRyzAC0hHXg4rfWbkp
mM7l2qW+GITpFq8214TLRSIOlvIegvw+MfPPTeHLVc30iWXJ0xv4XKMIF+cRHv67
RUJ8t8hyYJMVz5Lbq+mXnNFv00bEhtfcI1uQrk7oLev0b4xDtl7Nrck4qT9tXNPA
mj9ohcQYThTjnZ1daSw/y9V1x1kNgSfKnq1AfCneA0iMRTIrv41IiVxYJBEcOos7
xsUI44pLPx8fmhr272kptt2Ir/EioXNDZbxFKff8UmUfkCgOzt5X4hJjFyX58fys
brPQRRc45C1IOiydQ5qJNQKFuQTC5gwDfZ7OtwnTsJBCyW1l8mzV/2J3mcDQtP3P
j02qH2EZx+nkBCwFsdC4fiITQXhK//Hyiy65C7dRBEi1uikT8t6nSU9YSeuRyhSe
gELIkOtiA+f5FjrhN0HlYYkASiXb6WTEbtAK4G1iajtOypjff5XLqbG6g+LxIunS
aJOvttxocSGrQzWTSgZnXMjhjnQeGhkeenf08WuiSySPo1y5AIRrPstoSMLmXbF7
xk6VFqeARL5gBSN7KQvVBvTHlGVADjKNd+tG5h1QZJQGhD0zvNamZ2JIutfu54nC
KW98O8tVf2Hy0Zdw0KGzmbgfnVmk2KMLGoiggfbV8yADGiJqSHe5NFeImSHwLDdl
+vyIx7whOZpiIYCE6pnMnqDVWB88L2rv4trWyM+8WK6QNfoLfVBlKiRcFbj8B7Ek
8NTuhrF1N7PCLN0j8er7F3ZKYXvCP/OGH1mdkmZIaBNy9t/4xCdqet02yDtdtAHk
HRTICWUhMg0MDQT+IL1bnIda+oBtyfPGfOQvjd0XIFadPEmXppTuXemDCu5Tz6yb
glWfeLVbjXuqVESEu7QS8kHEtJRfvrVFJWiFmYCkErAVrCq2H4aZNHGw/5QTvrB+
jbB+xKhHLMz1iIWRafcyWA==
`pragma protect end_protected

//pragma protect end

// synopsys translate_off
`timescale 1 ns / 1 ps													
// synopsys translate_on

module `IP_MODULE_NAME(efx_asyncreg) #(
    parameter ASYNC_STAGE = 2,
    parameter WIDTH = 4,
    parameter ACTIVE_LOW = 1, // 0 - Active high reset, 1 - Active low reset
    parameter RST_VALUE = 0,
    parameter OFF_ASSERTION = 0 // 1 = Turn off PULSE_WIDTH_CHK assertion for a particular instance 
) (
    input  wire             clk,
    input  wire             reset_n,
    input  wire [WIDTH-1:0] d_i,
    output wire [WIDTH-1:0] d_o
);











`pragma protect begin_protected
`pragma protect version = 1
`pragma protect author = "author-a" , author_info = "author-a-details"
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.4"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
n9GXfY6k/ZhtJD9kiUNVLtaH0OSdANAy0snKnBtVVWQ6QOE+Ndo/VTZDI+hGg8g9
BQuVUO9VYpfcYCQvBCADNQKgSAqxFZjzIRV27HIOeZCFcQqQWxv7S+5zWngR1OAV
+Gybs11Q3LoZ/IBIGBpd0XnkdyubJyu4oBd3pKxGDxxRxImpbWTGclPoIrWLQbHy
BHYzpKNiI06B7YEvoi3X/d1pKZDVylZEMUSddSlug+uFiiaJtWQh6NA+z/owDEDE
V6bVUxyNm5aGjXjEzEECUcMJcfeV956Wj1jl3fVxGiNP0REOhvPr0bI/Girb6uQV
p+McpZkCfrqzEUBv+tF25w==
`pragma protect key_keyowner = "Cadence Design Systems." , key_keyname = "CDS_RSA_KEY_VER_2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ANz2D8YrxkPjLNtSoqQ0qL/n/jE0iquIWk/3e3vE+oIaj29rVvK4slX1wAMRUX9N
upY9Ha7G82YH6HOWpzJQwnJ2DAY0Z3VQ3OFLkDk/Huz3SCQACFeCg8JTJ+gkqyIY
3qkzAdDWdipMtrWdFBeESV7jsaxlunckrpbgbEzci0JaAN21i098RIWuzrZr1HTH
dhLLzlbWTgr2KnB5l9x0HVdJAN9fzTDmnCmAJMU6tkoHiQaAhQNuBUDo0LAEd86e
FLJDJhF15fh4yrlIrzYr3WEqxNEjnYmgMEPuSLo8lQrcsVIomt1zamkCO09pKhfp
/GUCfdkRxv3JWfTNRFn7gg==
`pragma protect key_keyowner = "Synopsys" , key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`pragma protect key_block
Zr7q0eHhaH7ptNB2EeBR/IQwCwGbZ8h5GSZSb4880yuCpqV3mF4LyVsWhgP/s+oL
K0Ls94YLsw+5IXRtW0LZarLJwXt3vd7exEKa2b4yrwhA3xkg4lvSFlzHYvUrejVb
pvELZpNMkl7gKvWAY1rITa8iFy4DIl/v0EZIF0sNnts=
`pragma protect key_keyowner = "Aldec" , key_keyname = "ALDEC15_001"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FuzzgfHyzdkm19HzCmIN77AO/gXQ89jPquRQ3E29Wuyahb8Rb3IaHBb2xF+ucNQz
iriPZJpxHjpFDU1ldMRZs9rmKQ1IEUkfM7Uriu9aXykiHujm16In9i6+P1J+GMdX
fZceSO0vZqr7OJB+4FbDAMjM/QN925xh5XTjFn6MNb2q2yn29Q7L3rCuZPQrb4Vn
lEQirmTxGZ1E+vr3rJPjXwz6dreTQb/ZBO4iFjveuPzjMlqJPyzHguB1VpgxGTPN
IqMyha9gI2WVCxiYdOnU3qGdds73SXmLkRRdn+veAxtnq3kfDb9Dkm0Mba9yro3D
hqg+l7kOuLXNiFKheBoksg==
`pragma protect key_keyowner = "Siemens" , key_keyname = "SIEMENS-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Nfof9ZZHl85LF7VV8kwqITImnG3WEZ0P0YVzEeGvnS0PevbCKwpIf9HZIn40pDjp
6C7dsnYUSjkFk098OQT3cxa3sB4nEQ7tjghscEBIcr11fLIYDU+4+loBl7+vKhSE
JRtG25f4RN7VbiA9wVAQvgQi4ruRsPHC7WogI4wtvEQU35OHjmeDHS3L+Wnepjea
LnfRJMDlzCoG/Czx+a+eVXCSIDfoPGZ86v2+jnHyFeDiO0Vs+tyViM9ODIUyuDce
hi1T1CYfxnmsbjBWvmVUO1sVbRzXnMCK18kgayk/a+4zZuMsazRunqrSBabjCfrv
HMYPUZ4HGf4jWmz1yLuexA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4288 )
`pragma protect data_block
X97EA9rZmQyVSKGVAPf+pA8CK1o3C81qFxKfRs0qOQR2zH+ydX+N77GBC70b5jxR
f7gLzUE4q3PYwrjcJL7/afdvqh0Pp8v/SNilbMnD34mjydvwzGjQnDJWuka/jhPI
e5SADgvXe1boC3wo60+VEEbdvzgim3hjcA7hVhnxhD9adPktzNj0IbHZc6g6XEjk
hXbjsrqbLt9QQ9jTpFY0Sl2YQIUhmZIYbwdXZoIOAbx+Wo1WN1+7JrB8skeHjcBB
Zhp7ZxC6R4Ve9wLCBQ0Y1kXORFPBVAr3H+vA3NSfCUkNDxKTkwsWABvMmENIzfep
mxUjjhSKIBBAaOMFFzqczgu1TP62P2uqtbbmtVZc3IGUnNNm7gb8E5XDEMDK2tuM
4AWtjwUpVVik/i7gAOI3zFboS7l4Ang4YE9oimWH5Ag1IF8fkh8ebM8Gm+TqGoRV
W08t9OJ/kps369wuNrvE8wTvDmIkVWmd4pLEjSmrEjKDAcsK2dAwma+u+crNEang
Kkv1I0e8lbMp9YU+d5rjgEE3czA+69AZMW85A0WDYUtBNzVWY59ipJkXCLGt3/B2
m+5vFKdGvN9BdYF0tFZl9WIbdYfNfpWz/yLkzD9HZDVCMj1/4rC+Z7smZ3zAH4Iz
ejonoDqTaJdLJtvDaizMubBK56t1dfRaFNo1lOI13oBCnmi2ol/rYegDtxhJtDdJ
oYCHI1QUNhv7zPXOIvbNdJLs78g9N6ZxNd7MA/7u/3LkSyXUErR1srif3lOHjK+x
yNqmvxxQ7Wx4qw4vs5/L2DVtHsR9xNjLiBs+7sfPeF1E7lmEEMuzoifMdZztZjlR
vH/bDoaTW66nJcERzXcX0YzMX2vY1emTeSUzAoqcFDh89Z8kh2OJLssqkTctOWT8
mZxiZQvy2H5iyEAStPYAxYpCe3K3Q6ht0sleCnJ2d1aWK+5NCSaepAEzszlJ3P09
bUKklikIflTi+qm3X+Q4AONTsKoggFCRUXHM6uOIA1sunoMdQhL/pGcXvGovEMgh
R7dve5fUyEA00sQPmmO6lJ2eolbCMj5vHqJIefTF+gz678wUjpkJIwg5oZJwktRB
IvcsT+/vrSZCtCgjOZvfWvhSQPSSfdws/u48zZ5d8nfhoKxwTNWfzR0BlPVDyfQl
ekxne2nwD1UxEANWbbXjc+TwjAZws/QWd9stHGdzlE9RkS4B+8i+EibHfB8clN/A
jYtwsklGwOediy+mmKi0sq40l1ebb68WYSdVW6+ZfbMzBEij5e7Rbxbtu3M6sJOH
alqy+Fanh27H09T2xw3+vcmErU2F/FJS5qCaagg+OHaKhYgYIKhdwO8wF8R7L9t0
/74wl8MDZSvh07eXDkL3xaCqDPbtv9dAeaGdHvwnEKciDafXkdrboTAz7nPcR6LX
ip8VGFuAONSaTn8R+AZiG36ogZdhOL/KGPVHnx8FzwIJpYMxG2I4pC08giF1T7yO
nHMtA+JTjVQPnMCGZ0jkMICyVT+EI6wRsD53w4isYqve9jukUD9G4FmOR55AR9V8
z9b6iQoSoQcwlU1fzqanbFbMZ0f6Nqmud5N7xe2DLzIw0LxoGo2Mk60dZPNJQsQB
INQOdGVly5oSNgRQZzOVsJwqbQLTbkZtrIa8lv/PfXf0iPa6xnfpDbdwkNnt7Q+5
UFBDpPQXaKHKt/EiJz3B1uspdPe1xfAoxzUOgusx6Hkb0kd63lKC3N0jwETnMCUL
PBCHnDJGRZphGHTVE8ZqL5ixKhKi2nPdrKO4Zk5sCHEpR2eJUobipB9Pg+wI918s
Z2X4+XeaTmMyYbqUZW8Q0O391gL8QBlmI2bedJp0NwcgIjbenlc5qIs3CYlFo0QC
Pywv5rSXuXdDW4V9JPsgj+2zX8ciiM32d8zwloDodaOzBxp/et5Tkr7jMMNPA3Tl
6Tlz5iA8Zt4jQ+e+qc/KJzRmBa1gmCG7bymv5XIYtKKgKOgv1+byxIdLYCMZGhIG
7kq9ctIXUDco3wC8mG+xXBWE+osZIx2b6l7TteZa/Zk+r4XK1ikGo0ukN71wN5fx
E3W10XsFdVVV2fp2LneAJwUUniG7OTicH6VlEfMwJkFMEroA35BFiiTj8s/C53Ap
Mcw//CzsL22voXV46MhPjqWAlbWf9JB9RYgGhfFi8pVVI2tXmMrZbZntavcYCsrA
CnyteYSgnniIvfLGWAMi+y2KqusOLETAjbrZ8BdN3fioKcQEnR7Qe5ePQlLKD5VE
JusFOYxwc7uV5TAYk2UYAdJwY6MaMq7Btl4SYb+UsHJfMhTbwwHQ0zsIW2x46S4A
CfVI9WDX6PdzxPCnYA3JpiAGL1JIHMzBTi1/l5yCJrY0lzJRAtd/RJELxaDDLbkD
Yx4+l185g7ztYG84IFaxpqXvmSWDkD/5t9w4WIsB31I4FcOyTygmVE5vJUsi3u8N
nqfndnyJ9yPmcmIQobA0LJbgxXvJPQsfWUcL+kmzwtzK+FcaNPvQ8lkkar5zHKlz
5RCyd3TKySAnX4q5Zb9I8Lg7zfwClUA96Hx64uepwonXw3+fevJ27HMDyF4rEidg
VKKKsP3TYq6/a+6U/UgeJe9GYxqzCzt62S1kde1TprEdw431j8t/f0cvdMwhRwhQ
rkKWZdn3lgqAWTCLhDdBtIRRebDauNv92PclN8Y3Q3JRtCXF7pOJ2KBNG19oML59
i7z2LcMUi3JgWWZyiyOb0JGY0En1BZ197wJqVOPMesOMNc4AeD5IJBz3ZLORlzAz
Rq0By8iVOJ6Z62EeqhbBv2KyTj2P9q7IgQDN4pvV3pDP9vpNxVq9DW9IDKfTIEFk
n8g8tSXRWE60Z+va+09fdi6P1kh5+YFbqfp5FSqcw/o5T53GjPExWUTJBaRFsPnQ
6gF4Vrs92wNL5MmVED+ZzowDz1N2l+7mT1s29sLpfUnS5IE7A05FNubFXaZmIyCK
oJH2DXvC0QJjocHr0poe07Box1/6w8gKGstjDRjerdNwfnHusWaAvx4nZorl014+
uzfSsqu1qFpqiJbX+7fB0F3Lb4VsWNInLYVhdlpm5aXotLsTCT0KmnybcTMq4Vs2
DqZJz44VhuauSmbLT2Jq9FReUGwS+KKn4/JvLAYuHAO+DIyumkexkvFPT/pAfajk
o1DMEHsOZLjcid1mvhgGiU32xuW8wC2bf4xVuSHEURLf7UIK0jDX8T9BHA1xHdBB
fLtAEa+jVTc4QRfBZgFYp4sNBwrXsV9NAKHV8HXX/mjketCpFv+Gb6sqQb/FglxS
Yh9ApKF5n+VnRxqNAxjhoBIKRbxlc/5KQ7N6oD0APL3I9I6oocJ+RJSgEk9fpLWi
sSR+HS7ypXxXgxmA0gTbkgKIABNNwyhwVAF+HU9vohqANOEJNygP0rzVDJby4GVT
llaMRSBt/pmlhEQWbCxbdb6lWiLEZLqlz2T3+I0PZcytL9LMW3k7mHKOBSvsscH+
IJHl+0m0O9bfRFlLCTPBqlULLllnFBqyLL3/kbjWjPUwMXcnFT812Hd4d4TcVLZw
CgifH0Azmw5Ryr3UH6XXzxhKgQmClij2YA343z5bEDeeaX5JfyhieSuDxd6/dpC7
X7FxfPwWLX8+Epxwj+A3J4a7kuxIv8sTEkSxFSheaL7BQYQdIbCw3fFqt5gFIeMq
YhBGKo/HxhVrGQuyep5y0QkZmH0lOgEf7yv9bz0iqmyTzxO2MgeUiN3YCg/6o7DO
j8hTdftICEWV7jzRjeG6KPuj60MNySwH0qiKga/FVbHoCCgCnbCJCVHIJ3V6Tjli
ODasI7wvSBWfvOcVDvcQhtE5GfDS2175NHA4e5PS/R9nsRaChoQYJyuemqUEp75n
LvoEVvCuXx2hHeoiXGCJswKvi0Vg68bbl3H/VXKpkFfp8+eldgVjeKuASbynUICh
8qnv2SEq/JZ5NPsBxy95MAlhqCaAT90gn3xsHzOSaxa/D1FUDYANVKYwSGO9Kulz
XV06VXPx2G6YydPkmZUnn44BiFtQQE6sHTM79reOqOD+5/zImBk/qNaEvQVsVXfM
nttsF2vp+/HTHQ3CdM6PoLAdukOpzkDzNzuaj+mtHT6/6tfozYzvE8XV07UIQnG7
sW5kEH321LvAxuLxT0ItIdE/u/o5NRPUdIpt6BCW87wbOVY4FFuHrZmPfxvjR/cr
GY1wWkNjB697HkUILocXAKx8nJHB10keO1bRcM0yC1mFfssRdbrg1xLxrJoul2Yf
mkhiGQjApD7NAyYfIOzQgPwEDQH52h/VC1403QbDqYIUVlgycPg67P2qADS3ObbA
tDJYWCp9DJBF3Xs0vmetqFM67rxZGAUuhGMGRVcMpFmX7s1FVaVv/7Mr49POX9XK
mv9n9MK6S2rSErofHE/+9xsFLS43U5azSwTgPnMiPCWHeFc1SxQq2yJR9tqJPhPp
8i87HNvrD59PyT6VbT+5VZq51Bs7/t2gWDzFt+owA3oYYckdo3nN6bmYjxKKmHtp
mfmpkkYG2uLehgXvZT/gI5gF6sIRh8Mg5Otdcn8OyHTOq/Hn/ngbXEpbfX3qC8r9
S5XfDr20ZKfs6943PqhFEccWC6siCvFGs6lm6L4R3dYrXgXlz6Yb6MOgP30GHIYh
d5W0kT0MpAaXP+zkyz6DH4OIGCIwY5BdBVPhOfn/dOqhsnnmccZdfj6RVYXK+YIt
Rd4sQeaMgaAP4sBIk6sveA3wQMKv6bfJiH704yy5yZnpXw/ZZQOmSAkspV9fYYYQ
mv6Guobuxk+KdlDcQ+WK7jfKVgdAAhgbAyh5mtu3BxXMZ724Kf6WYwa4icQ7/83c
BUp44S+ljdSRYo7n4speThbeAlSlcGGMYoXaDPJcQHpzAVbcO+/JZu8Jwpews92x
wx44IY/hTBZZs1FL6eI1WoqxUH2IStzOLP7MgdkRIKdCUttNImaR2OyEV3CR37XW
zhRDrP4m3NMj2YxAvRqAyrmzpv/bfNmTIXbLWgeuCE2Nuo253KqMqaN0EBoVFs0T
QfivBCQhQFx5g83P7GZQROaQv6QzRfSyPfEd/OnsX9BufCjiOvTWEU4U1hsrr11S
pUrGDscFKXGQnlRkn9mhWp4eflCwDvdsy5k2E5EMV21opUS/wIybVQY5fQ7wp+as
8p1bLj5pC+pxDt+UVTbB1hKE261Hzzam5EeTcjb0A8jadAGZ9pycWUCNtF7UCBTX
Zaoz4bCQjroKB06VktHvDciBF29valOeuz08hVAls2ngSydrAcEBvXPwwwuKX9tR
bA5rRpM19xXDBUk5NEi8sh/vDyB8d3y3HcdQyEnlmOfDoloY5Z7h8oi3ilcJQcGJ
8cOzXarjODunJOVygKDyhZEca5EWEwDkx49TGcPAdE5Jnw39TL5cxac3ERxX6ojE
ZgR8kM6bBuzNVdcIQ/n6OpktOgcpoqb6R8Bz4iUb4zVBGFqkrYFGyzsbtVn9QtUa
jhSxj5FiynXJjlVsNNlL/1ZVA7mnXXoBX4cX2Fv8KDev6NLzqKPwYbiIz24eI9ya
1Z5TYyCuP/0EZLdPCNUZveNY4RspJFIQuhnOSIvPGDTJsS71I5beJCJ0bur01zDu
/Hzy41OwhFkW3GXBgwtgZqThTXp2t8BPdQfiRjZWFL/frfzCkCRdJkOY84Iyugm6
e+X3is4RzltxP3oHsgBfyBxTaMedsBhoQVW13478CX2kPGk3oQ+xUgfeKpwDH6mz
A1csd1tPOJMVvTV2UTAmlw==
`pragma protect end_protected
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
V/Jeo0iJE5h6sM/43GVwyL6E8HOH0fXUVkUie06C3q3GfP7WCBeo0J/bT6PUa/SF
66fKU4Pp5LPDwbefvee7we9yFdTmaOcotNf2ny2C+YeY8i5qT/BRrbORMac5nZSZ
1euVfGiLX4zFVKU/HnYFQpgr6fZ/mc9ZoD/bVqO6s17L4GLgxidAWq3+lnLLNKuS
FErxgBjkPfWc1v4f/vYRinwWsbA1t+YgfEeVMXiReY3Gl78W9Zf2hCtfZ2wcAe/c
9qVXIreWxjp2t1i9NpZQdQyRgdmtRL7Gcxn3sEsqJW3cb8+VpJSkW29tdiQfx0Lz
Tf/UC3ywjDG8oOgPBtcgmA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 37024 )
`pragma protect data_block
ePTBUOBD/oQOAZq7OXnUVoY3B5JKBHzquoFqdYUt37TtSSPW1RmihoSiWwdBnlpN
idC4UKsKcEzkd1zXwEfsJUYNYxjC+2E73ApS6Kpkh9oO3QbobdMJyLEMTX/KHTyQ
SQT7mByC6vHtg/OORz8btlf9U7aMQxtjX+NSY1JjSFOc03ELpvvdhOYeaFkViXfb
k2EzY9cctG5cRsByxNJrIkSHmzn9t/bi3y4aBx2MEv5lAWFZ2uz86xuVD+lIHDYP
qN4WKB8WN07Dse3MdxDw64+aO9ap8AY81LI4jkSsjcOGrzwYUrnFDzXh+k91VIgz
MAk70Ag0dlsdGs69JOEwUmrQrdP/DRBbek2sc9q0/bF51gpZ4dJFgItSCZweFqUV
aw1NrG2hPQrwmWCj7LKGbUA0nk0x+AOy88jh6G2vKMsJlZqHmFz1s+iAUgJgpssH
4RFhW6LyA9LCIxz9m7slumcIuSzXnOUdb6rNKyChNv/RB7/M8rkPMRg7YrtveU0R
vix4XElEnTKv/O/8XMgAh4HWYQnV9/phvee3WPQQIrfKV3b+Tf77/X6pNl46IspX
UsC8UsYz/LatKrsSYBtiQh66oteAV5KGPq35NnOvrrYhReg54eTeHMRXrH1WgVb2
zRRMOYZPrlC1CYtugh7V/w7ekgoNablkDamX4DCLnZPOVxIIYzTqdEqhnbHnR2pW
dQuOQrQh+YkBAx4PMTvqLQLqAqQVdLp8FH/oAb3yDXKzBppmddRUQI5n41ggHCXJ
9192FGlINlo67mOWOR1IiIJzsDAgV2T59rfEZAq1RddazulvjO5i452pOtTvztRx
Zo6TPyvD1Q0Pbkg9CJcgZ4Pb+X8y88AYwLHjmmekAjLj5n0EQ6NSe6X5qVEtS4Bl
1A/XJRRBMW0EmBL8RNme9FzAfPuOmj2WkGG02Rdmm66RYPlkiaq87hMIB8P1kXgs
q7lggFgovuVEeag5XbxfQaVojiL55tleAc/v+viqnhRlEjUuurpTgfyV2uePB0Nj
QH/F48GjKW81/o5BHooVGmERdAn/1g8bq3ssBTCHe4wRN8OaJijn2YyrY8eaojif
vraTfcZpoA1IjnvENKAa6ZwgMS/XdKZwj5nhI9qTHeUi39wDkXDoM3MALfBgWA9S
lOxGcmz9S29vwOwloH9ZL5fydtky2o/fbSQ7f1DzNhzT6TatotQAHwz7SHh3IPpd
WOl1WG3IQfFuWQO0cQOCD4FBrnr2aI4sC+tLSKl42cvaEGnmSYk9iXBDsPJYwfLb
Ju6imPk9QXEGHZj6TkQOLCr/4jw0n4VcXFS4wBNMw8MmT1m26pqadVMiN1uSgZN3
u7zKKEraBX6hqOuSgbww2H+DBhd0PBtDwSf4qbStAkdm6ilqwnQla29uJLSAEJgt
AO5fH4UALWPalDpW2QZ9CEqsoNr95OBGGvY0bHuxELKUNfYoS77Dbt9oqyz/AEJJ
dK1GoS65DZ6R4NUu8IrHjiT9+SMqlyxwrqR0QdP67a7IeJq7Wukvcj6J7JxEcfsR
41gnEcT9BT4rzBKc6mdld6VBhFfHDSqi6QUodPT6vEM0h4Gsvo59A3SunRC1Rx/N
J8EW3O1paRtMgo/FCBYJ57QITGEMsdWUPLKzbzyVQYk3QKMAR7GUwDLKn5PmzrI4
z1Nrwvq0yuEDrPf3d52B5IAlYiPnViolD0Bimygd9xbhzkbOF6MJi5bMWOJNZNHP
r7A+5lKu7JTR8lUSkmUEAYDSN/1h/WyQjHyM1SCTDX159PWaGs+nsZV2gqTNaJgq
s6BYaLsXzcBqfDfeVNV6qrxLXYVR42AoT6D5GOw2fZEqzdMab0VXXwAko5fDiZ/V
rsPuCoQyK8NKq327QA+BE2X4GSHNw5stiCmuYFSzkDlbdkpZGyk93Lmw/EU9N+uk
59VWEENSkbNwcCXBMnjAm6KtvjmMZ5xffHAlE/g9OtE8t9AGG2K2q3pFZ+VP4mcu
ll/jyOgf8bqp6nwF02czrKBAG1rUnztUYxrn3ezV3QqfYf4wBaJuNMaYMYfjjY5f
wBcyElb1M58J77qiJ3wZ0td79U8BvjidXdHedxLw4wgzNIOoXtYiCkKVgTMP8hOE
hfnW62v8yEJnAS1vnDPDUrm5+dCKSpXlJSvFae3U8+YejIgprA/bMWY/OcoXyEAa
WiCf7c98rv281JUV81zjYWQ/z6M4sjQBz8aQbUArFbhVbAFwuo4s+bOZfjfSB4QB
+SevRZ05VcA1hOuWvkTdhu8LeQHXQae46/ocxxxDy/qWLjEx1LAvGL8levFN8hjt
E53oA+jaNdFnMWUq4Q2g7rRmkjc+evfCBM7Tw/XhUGM+Y7rpaVO5hXB1jLO5WtLZ
qN/L8GeKLTMdSBXigBZn4s8pbTKpWCnJQp36OvPwmRSXkUC44FEWZHDMlI9ptkw4
LsjWL6S20ZXXBJDAZ3w3Oq2El3RFywqjzuNH1TBBOISnkBNi3v+eEbE3Wwqy4fhR
VOJdw6mWmGDVa7qTIM4n2kS5IlayAE6hzy0okgZUnH6Fv3W5m5fYbd4+mFkcomF3
RTuK4atvwL60aU+8klIXdkn/ARgkTkv/yF9yNhGJUXQvvCscXmvKZTnNTZ5Z+066
RbueMfgQ58r8bEKi3xqDQ3LUviIDlyysPfo9V5g6/SprGbnRZYpmYhC+VUb0I+ep
lURY1eCawElDxVyW+RQG1ZbyheNum0ZtAXMnVPq2w6dduf/UvdJyFybCucNaMca+
uJU8wSPw6x2W3p2dTo7TkkZrCM4fkM9gHiFl3tN6xuHrR8XHz67VvP8FWDKK0uot
e+pjBbllrDUgxjrbmiLJBrhGfMX3y2gke1sLVt2iA3lGj+B2QbfWDpaJUOLbt24e
M3O4ZF4ywfUsCCTCtsxfO+Uz7w98G736sAv9QecRcikgYxXGADBF/u08xVLpBZeC
oZxHZOil7WpLwlKHaHeOTaHaWFVasqT8BqKEbj41Lnjd9i6AJVXC+H53DeSJnLjZ
YzhJJhvkkE8MX86B4E1uxyb9c2ZMUF03ZWs/jca6bAaX3ABa1Pmll/5pTvwDcxjL
jwa5tGV9gdEJ0rR7kU8O6HHlOSr9LNOx3wX8AW8MUa1Tg60HIWn6foE69QsMqVti
pmniBG9kelobFZXzrCt7On7TYmLrZcyJyPB4gwPz08zaNXDdpvG0WEHmA1W0zXtz
NkJDCw+ciCl/QuExBow/AH8UkNDsHyE694VVI9RJBJ8JwMn3ljxIOlTT6AGqzChJ
5JKQnTi64/Lt7+2OcLo0PjxoqcTV2BX3efdyeVBLQkhHIxrAyFs6NzZg8GKw8ODO
/dUkVtZjO8DnVuq8r4VtAm+RVmiwMjrSnMhAzaBXoD+8JJybrvxPuKnc4mg0sh9Q
AfUMz94dwWe6io0YG7SmGZMburgROjJ+D3K8baLRftPQrSUEDygK5WASn9weWVks
aj7TBA3nSXnFKG6NH0NvgZtt8SbHA//fISIJTyLGJQpRZ3LJXWRysdMxlduhjEFJ
voas607ZFTjinmGWPxgZPOok8CAgzz7OBSeYuLfnXaIw8/TELDk6Bcc+aOn7V5zv
NkPSb/bn9I3X4rYIxaIRyAD4ZURsEwse01NXUi+O3jE8dvipitCSYf93XK/tLou7
+ZZDu/w8OrbHa5sD9mQxgX2RVA2Gcka1V42liBvyHiNmEPU3WMsXF5sBdTB/Y/UV
jJpIwUFVnT7pJIF6uSblJcCECqNHKfx/NkMkEZQZGDIT2/v86gEMD99G/Mx069th
TtAe1P581x4/oace1CFZkIP4iIZwywrD3lOkTHA0qGkkaMVGFWKMfR+4Sdl3ACX6
o7AdcTm5CElJn4PjRh6xbwgJjgz1UOdDtdw/gG6A0QccM4+YmVyJ8awmNJEqLTkv
4j6N/I6w/HNyrAlxtWz85iH7MWlMNMBtnJBLXA8DDylVCLBfVHpPyl/p+wVc7/IT
U5G09Cr59nj+Pi6wn+KHogtwEByklAI8v203tZzVxdA4nP4ddixu33dUc4uuiEN/
3VbZF2g4Cki7049wRYatZoqTNEZgfAm6/6JAYS6Kmoa5cjsF4uk06XuIooTiXrEo
xMb6SPl8S9GJiyYT57mwrnEEr9n1H+gkQFgrllX81Io5UpaoK0yeoedJuIaZ7nV8
wMNpIsOI1ACmMdJ7u+78wZaNxMFd98EvbMEmctZA2r0c6HJoQnRTISVqJ1+2Of9d
B3FNI/RL6/AZx1Wp632XOdFpnIzrqaHpNhFmUfrU7ukNEQNwOovB95Tuzxgcu7BM
D7qZ56LVGeLhTDE87JLactYYr1smNPdPwqtgLyOlhb/4dfzLZs4Z3cjBruFAQcSK
0tuXCTMVm6LBhvYCWKD5C739jAiezRBKJ1dXw0V+6Al8jGsmGsIUlWSdqQiO/gzm
ecvwHrBdSoE3wGhRzj8sKNjI/fw2gmf12huwhen6+O79ZvsXEbubmEBdC5t3ZCqk
UWupJYMugHWjpwqR8nkojnzWVcPB+oogJ8wMWrMKkhtkrlUHDC+L/UNO3HEbc+sB
m6GIbFnhulFQLFGYGaayQbIS0eTkcOSQwwqjVDC5L/f1CsSkGIMDULb4Vjxstkkx
el4WvpYFP2ZQpR8Kaith1J1Btvich8gut60lp9bUBHbukoR3I7KF/RZz2Z89D5Ei
uvb4UNDAxcKAZvUypaxdW0vTzhqtdwxX+jvD4GacbUCftdJl9mtDzpwRLeWTYpFs
hSQNRsBAuC+NG/FhZjiTTgzoR6MtGqmeYaFoASE4vm+KYxbacFAT8zR8PZ7l0HxA
8tgyNg3VULnoSVheri7adLfSkJ/bmf9ELFkOKTOQy3QpioGI1rXtgF6Pz0fNw84V
XLElJo9PgA5dmpOAG9gPz5DtTPI4iHz4lA+DcKEu+nQ4XWRn9u3bRmQkBlpE7qKa
5e1rq9g1dRRFdZ3K9wQT3JdcsHgOw/e+VYSFWUZxSe7Djxqklk0lueAk2BJhB18Y
Vd0R1MBVm5VL72ldWsHebMBIUvO+VnmHVUuF9Ebh3QZOHr2+LpChiSw2FtjGcvj6
uYnwZE2KFAeX4zQQMzPUYv5Es31srYGxa4Xn2EPc/tIEkI4ixBvYB710Qa3Py4oF
tDYIpMxQo8unRJakUQE8FSzZazuiyOSwWA9fnykRx6dhHiB6N/1c8GdSmhQAlXAm
VmWP8RMxYeLQAYAHQwXQ2w/p/lamU3ZLwtwJKMZGPi4nMOtwAJ+ko+6rhpulLLzX
jcNpsVKV+pdO6veExq6UaRv9or3fgpgdWeouLuiDlKgkgYv06BRjlyqGkFvgxwRP
pfruBzKB/Sd0VnS4uC0Q2SBlaWT4k+mb/YmnJCXGZMS6jX/fNqAHlCaM0PcPXZrc
fXxZehsfVUYoPA8LUrRgZ+Rejept6qinSaYSYCXaWCWuG7LRLaTFR2UQGuJEfizu
SorAZrogoJw0Un50m9I29b/Hl6zJpf8JYF3SaKtbTGJgvCubw+U3y8AIG5ANZtv+
XD+k979PWL5SUr0jqkODoj1jtcV+g+8n/DBEaPDyQWXqKLjGsEpVOphIb8ZSo6LQ
OtX8/hM9e32l14yqyOLrlrsbVwAs1VmJMvd82w2vpobNCdGL6jO+eAXF1s1VkS+o
1njQ5PMvLWbd+luNxsNTRHCtQUFwRcvoEVuXRnQG0GABpRZxNhFlS+ia5VNXAWWY
yAWJqDuFxGM9dCLPCI0OSD4UYVOXhLgxY/6vvpmxt0HyS4/zIWGS5EU9LvIbtA7l
+7HeTmVPkigViYF8dj1C8OklA7JEBJq61g8cYh02jXskkf/nm6bk1k/JwoaxWQh8
CG5jGl1fP5Rmpz2HGTRV+O/w9SQCphZ6i6i0Z4IU/8Y5+1U8QWntEPhkvnLWWSo4
Gpz/CrN2TAOEAaM6frrdoVjZXnJd7PZdB8VCrluP9Io59qB8aG4F+X2mK7+aN0F3
tE+PvfNBASb5o9SeOpzj71vOXE+22aqRG97ALS+r60W4fYx2hWtGXozZYRfw5xBs
uHXP7uaa6iSiKn146iMHZWAVT4iR/YN9SSNy2IH5V79RL/5yXHQRA/4kn9QDVq1B
zJPU6Ww3F1PcryMShqcbRwU5sb9OdHNJiRrTWJCK/cAPYwJtkJMvrh2NwIh8TfGm
Pbl5N8hfnvouAih8dkGmif88DHy03BtCXIarGTjJfDtg8M9EG1bOLldlmod4OWMx
5SXKXt7OIk2lDj71KwvBiGoZLDKmuDUrIoq2OJ8GF7E7k7Fd1LuvHbeQowbWpp02
/RVCWBqZaWOj4LtOx+xyrbVVd7AKwU4kNgMGstU/pu1ps+em35JXhN7PRyzLYxm0
KoIwj4HWAMglxLTpYJqdCJvspd5nS4qaVPFvfb5TCBZ1EI6LPxw6FgYdFPX4z5yb
wnitp1mqzFJH16IGiAnmnO5DNDpFCsAwJlsQLw84EhWpHRsmh+1qSfHuV8gKDE2P
58/7ZcOZdLHdVyqc8nlc3d45eMblTtV7kzrCCVR/n4VrD5hkw8UlL3hmDm5vg4/F
xy96VHPzwhkSv6ZXeYWoozRg6x/9KI0090ADVT8O3YoarL+4EthMYHPnZya3lKUS
b+uRVVxIfwaYHkqMmTPWyzio60OfAKzB8UgUg3VrCxr/dctw/4s2MxAldkNJc5u6
JLpjQdO3G8bjMXPPq1e0Nz4eQqfBOiL9bwOGPggqRzDYLapzUTcFGqKUJGC4Dxc6
zD7cx2nuXhszCYs+AZDx6XEgCNb8KckXem92zAYcaW8aeRNG8RM6DnqAjySufcXd
sLIVUjs1lUGoOX3u4DuvHvVZABTPT60GMzrsmuDfLLBupywmEG+nhzurB/v4YXov
v3JdwyVraodyyNLK1+WdmtpZ23q++1KqUAKtGXVs0AWd9K2/hfQ4n7FUIt8FJNK4
2n1IPbzYD5MARoCuZrjBmeDy7KPqD+yDejIuZr03liIvK7G62UvHkvn1Wj4zJdYH
R0qEaUC8YFXdCHsBMzA3ZsEnLFkux5C6TB5x++UZSoZvsqmND6t2l/QQ6eyE5Syx
yI9qTZRFJvOWDY6HtKf4UmEAOOnhv9O+w3Bk77TTBcLFNe1AOatczHMN+wPx/jVI
kOW32Fjj1fNxpFJUUb05Nwci+XTCdAoFh2mYZTFKLsNaUOd9bho5mtLf/ldQfXAL
7xeBiDi4v+uJ3Mev7cSU+vxHaWkV2K0CLSMCyVAV+fxnYa8CImKIajC/titUL3TX
Fo9C6oxDKryS9gDFQaGiZZnbmGKY5ltMJVc+TjV4abQTgAW31Mq5ahzqm7MJZNHX
rEneArg6waHIwQhbzqQaEq6o8EcvsUFcA4FQzJaP7TpxGKZy+y0WycgZODAJ0bAN
WIkVvnAFPrnWmK/oNlZkQumYcaSYt8I+RuD9ij39hsXmkAt3YxGJY0Zy1q/LpFv0
ZkH3iBCZkUTrRSfsn+InjsNRq45YgSgO+5s1yakuWbqvXt6wgwCwaLzqTUvw/GLq
CapPcq4W1Bs6e9pluW8MZL5KHWJzH7nyj1CpiQfRhZKNiQxFq8zmkg/OfBejOHsV
Eo7WPTuAgJS/qM7S5tfqQa+c0t1nAYfbbZ885NXEVVIqshGoPHTEpKmxCwoKu1o5
A5kFbCv7342KmtQTVLpspnmethYkDT1dPiyeCjmCI/EBxJd2Z31duV0WCv3pkcVo
qJwZYWeD47+R7ZNpkjcmeLpsX7Dqas3f7aS7tsEC8ez0eIgH2lm1I4exgddqknBW
wDyP10QNPhmc9Ym5sHHngjcxW7od9SkbUHMUWp6FfiLWA3nxwiCX60ze1spw6+v+
arhn2oayGGoWhfauEZeUPYf/19s4SOunZf2QZrUc1hWjfEABC1WERVc0wmzs1jp5
mj5lYS50JHxG5UsatzNOIUdqIx1mG4tRyzZAh/ZnboSLT2gmvp8i6a0P4vNC29Db
gLXA00eKgwAZjLEFOH0cPKhnJmgjl7fFWBAqJTfrOY8+SyGWuikBGcPBMoPphQvu
0e0LdyWGEn58arrCrXv08v249q9QqNiGjAdvyztNtYxb+joVI7upjI8VpaNoI6//
4toN1kjoC4hqlpU91g63hKFS2Zwk9olDnjbXXDcbhUijUsUHgQ6Gk4a37jClZBh2
tFxRh2mdx4BjLHi6pqGcoh6ud4PW3BFjP0W/UyXVIh5K6/bQ4Mb2eKQv4/BhP5ZQ
fbIDjOHF+pfjMQGzaevolnDGxh+hMcbvGMM9Nzr3nWqZ1UyfG/H9IhM1//G3gnYh
Sj899u2/1MhD8UMstJFtO1rNKr1aHr9EG9XlFXhKnGuBQdGsOATQcfxSSIRO202j
kYtzBZnOPgX5agXBNjzxg47WBCRKMz3+66U5pMFEdrV3obPsExAuWCGg0ExXXGTK
QuPYaBwI4f9q2HnYzeUCa/6QivvKLy4S4VoZl+oMYhgXnlTEBkS6Pa/CKwvRrxCz
EjjxpTgWbHDRm1rZOiAo/jzAslQMj//zhOuoFI7Qpi5Ex+fKahlGgzM0yObPXwwq
utkDDpx6jFrlOhOcYRDxLqT6GFf1No1cEL8d0M6nMls31BsFLP4zDyLluGUCdOuH
zR6GJzrFiBiTvX8D9vB39Lu8DgUvr/JkPD/f51GZrh+o7pVFPOZHhqNmYAN8ki0o
awRmUL8tzXcqahEJboMrTGfVAa2MoE08a81sxPKp8pHwyo8AkIG7iOnHvFZOGL7f
i4dxRRZLxtS5UXDxwOW63HEXKCCafgRPNJffYijt1cP0sDgDRaZUUkk3u/8GzQpV
j/jGYAhn6Urbm9iKfEaOT0pBYBBkzsjcnPL7CGqggq2UkLR2sUDUp+fkrxYp6Azl
86DU2ZRb9J5F9aGkDv/9VVkobpikiJn4aWYmIHQsZJg3eFuSlREnsT1ciwmEilhg
rKFjfSSLlM/RrjOC238XD8uq/flIHlUPefUM/K+7CPPrcY7zOSq6hXK8WvPl+3Zn
BHD+ys39gvXOcDdh+Q4knapG2xRYVkfLaW6zPtOsoZlnW2OmISHkTcX0NA8P5Fd6
NHaXvuZBE7uy97TXoeHhQAqp4J5REj04oRmPk1LgTkP/4tt60ma+SiALaAKyBjXK
ZEXuszQp7mhM8tXQ+pzT+JF1EzZY8gR0YCfQx2SAIb51Nz3220+l5CB2zRN9zxp3
WCUXnJHbpeQQDJw6WAQ0klHh0q+6JXGi9Hdt1DmNOlykD5mP09OGa12FCtfYWc/6
q+VqxBNUSECfKvI2abMTFW9zetUWxK3KAFZgPrtphdxQXVDM0Fd5D/s8jCGlrJyt
HJkM/wrCjUwkdpBzCUvIL7h82s9BCg3LGjViotoPA0DECbgGUYlFIoek9kGGTNed
WpQqR9IijwXpfoV7Lx/cGz2KnoX3q5S8kD/obfHVS3QsNefq2vvc3XqCgUrZfLzE
ugS9JB2qUaU6AGkXlidzmfBIbvO3r6nupb2444cU4E+ea/gqYi0wdFHQA8rw+JmA
Ve4CXwwKid1yASegaFtMw7/9iOyz20MjOwvYHWpaPgDw6n1Us0WyX48gTSTJmzAp
FRWyVBEMuky67Tqe/rpPAQOwAC3/1orwlNyN69VQjVD1soewUE+CGFQufMazHuuc
AmonBwCxh6yL+9vuiEyczkXr4fS3C8l22SBIlAVBdLs2Hh+ihOpCLoEarku0cmuo
DCVbaCDkpJfMYdvODezLDAjP6RlRy3AZ7dEEQbObhV63oVhsE86Kqt3KrJaoe9Vs
aXm/2grIiZr+EtMclSyJSK7iXYBVgXtchC76bWFUFRG64oZ6F7zfFrzYXFUpOHuo
Pyb62JZvhTLnEOhb397c84RjyThSvNi+56xSLb4XORGrJ3AWAwQPU+nxgRwmDTC1
JbhcS3jeZdKJyB2AaeDQEMnmvKM0KUfC/n2EYrbyUA1wcUNXMojPXfkh8P6fnM3j
ljaRdFxiUtP5IzkHAw4J8OkiIkx/MwQpDE+LwqfHi8vB8v4eo4On4vZDlpIsb/hQ
FVruMRsqjMNeufyp0gw+g3nvOnMk+tY2cxVznv3Ar/YE9UXuMUNeeCiUXP9XuVmx
gnxHPU1pTvKBznDTabeLZR4gfxvLmZTysvEGSHH2FRp2poa4lLodZcSBqUolDSsY
OVs+tQAW682jLB+Gw5Bl2xP4152OAvBGv6fUDsPrqdy4kI3CL2Pb0WQp3QpxgNsb
TyYAGhf0VAyHwTovXZbhw1DWGbt1Rx2RW3j5vQ+XNhM9VcQrhf14NaFJYHGOKKmn
eOd4Olo1gGo8QaVm1uF0CdvQgQQFCla7pAKh6u0CHwpx+NmJYP3icvCaPmQAyKJW
6EGilC9xwIkVDzBJoF8APg6BHGLQeXbw5N1F96B9qExRFza0BHSD+7HN9n5DXsRd
woDcI3uaztGvHwVqEBUgpzvgapQPYFF41JwYLLHgjpPYCwznpZNk/RluPo1VrKtL
uydsKDE9EkslYhJmY5IsSWEf8o4QM1r2ojv8g07SgVtLTcnhSfRsMN+4nMdzhxdJ
O4l0jJPWCnqrMcbq5PajWrig90v1UsU7hk+xUJ+ZF7Pc0DTd+ykdvRNjkny2WdRE
xnJTwqongIM8cFU1pgHM5jwKxb1q9wXFiEgQuGNrQ9N6nMWAOb5vRIkL1VwsNSAI
Y4hQlXt/AUT10gStFPt/RunVbPhVtXoOdoZ2aJEw0JegNqKDqLr6GPd0GkojfCju
ml0E9lXanyV6Jp9G8MkgZfaeFW9BjjzIVHwoJyxaigWt9z92/x2imocy49bdSxzv
M/VokqtfNjRVkCATtZLjhMqxSDNAi22cGN8eoLNb8qrfQ79lUufVxlSK8d6EzY0F
0WC7uBljMZaMqm0l8VXUhwd2l8nKhxFO0jm6VhHIbmvB08x5J00WXXwHWV30V3oV
8MNp3I1NAc8I/e9bbEz4ivBrSCILJkkVxRBqJl7CgfFpTkFnvSbXenZgIy9fGx3u
jXX1kkmekxIh/mDopyc1OmpUbZNuC35zYqpDEReSbnR0yWkX68ZPOAqC0VrtTBU9
P1ZmOzUMdOlqnNuIjuyHtbiPn3jnBDENw/sdlD/eYqb8bc+l+nIO/kovgXb8TsM5
NmhbGHrD2jaD/U1qfwD4rqGvhiYZcuKXA71uggPNl4qjigfakLDY1s4vYSx06wVT
Hc9feyVWB/wkkzEE8DzkLsuJYuRzaZfME1sT7rcUVSEqF5sq6/bgix/22QCRlgA6
wBvsZEwhpQ1FtoyC8+wghO7RIKnxNoTBfJ3dL9P9z5LoSJ8kw7m07FqPxcbX2A6k
GrewXKHToAJPGsinfubKmSxgLbFYyl9eOr9e4DkwfakZH3R4rZu8S4NGm5b/+YY2
QojfjrcmQjKvSqcqY6WE4/2CCnk3AAghnP+J8N61j5CSoGupMroMZJ+xZQ0RFaSt
ta4evzkqlNSHiEBxMc5VPJ9yiQ5FiYijuLH6677+LE/YHL+nCgRpQ3X/sFlWmYc4
GOJimyAXCxNENbHGXFNwh5KWGzRIVZV7gMYgWCaL6bpDgMwxpZx6Eo/UzNa+8YQC
+KiTMH019j5a+VvoziO8tmrMAF4IlWlwfueHE8Y7nZ8escLsizAtu9T+bIklo0E4
neRAtlgSHRyGgw6Bgp+7fTOvpYOlDISj7GbpI4HTLEL3MvUSVVhNNmfROqOztRLj
yeIs7UDK0elX6VwRjRLpZQNXSJRYSdxgEJRmPDSgq8KEfcgfDGWnANbs5qAbEent
zRXdGoCSKIr7HJs9cBnDcIDR3njxeW8iJi5cae04+6YLliu8jJduyf+r22LJEDjI
w8gTq9rzWmiZxn+k6UVErVjm31z+z6hMfxRxdjh730Q+NmEVm7ljyHG3Ahi760sD
cCaPbhE6Qw7iBEQEjJLXwlYioZIsR7Yl0w35/wAmranz4MF/lhV1K5Kjav1Fs+7/
EanQqxkt5VZLgMRbOvyuo7BlpvHZH3/+q3fipRPXhf8oYiL5mRZ/5mj9y7qoC/Zr
5fNdJUQEdC0wmVU+Yyu4qX++MdopJNOtv5y6datMHcfn2ULBb7AxTvPy8/l6chjF
f422AYs4K/62dFIOf6/bUVOd1U5Ls/glE+n5oWEXAIQbLDyeMK63avgiVLx6X+W9
4iOfNxHbb9VybaIVjIWPqSkcFEAOKp+r675ORAsLv3pe+tiupIONppQsFeDpcPSt
B9kPlzW+R19+DBBDnCn8tpiO7gLosCl4Y2Z9ppFn5YYnVy5g8bfr29za4m8xrU3s
pqa9WZFE9etdeSIVh+4smL+Uu6VkqnPLvWMLl/Bbssm7TEzrOS8ObBJfE/0WX9zc
O5pCqQ4E4WtiKyf25QcRFjiBbqRXkjKJEHcsun/dem4ReA+eob1n1bTSmJTMXtVC
1U1yUYm1eZdsM96Yc+90YSg33HkeTYpLnJUnp6ge8/+jjqcmoH/U38xszYlRgR/i
zoWZ8xpJ/g4RZguYcV+pu+5jPSfy0dgJ7WDdswLcFju1pzFy3aTJh3X0Ex6K0Apk
6bormLPVUrQkCFoH14w65i3hirSKtMb/JfPsCk1UNYPI7m582hNimj5u3yCXvIsM
BZjJajnWjMMoaNQCYrmiPTtCXqcTBl5pAFGAVa+1YKachk7YqE/fQ0rY5Tmgp6EI
HGR88ZeVg0M/x6CTi/g8IK/SqNCkwj47QCGIDhlWJU4/RqQPZOpNV6OtMYUkpWRk
jrXw7b15MbmqCqyZWLRX0nss+63TbaCL5t72JmwvdvwoTPEAK/aDm1cdpK6gtawy
SHDmaEqguIeLf8OvmMqsMBIw9RsCQpC8Ad6/6cX7l1ekR80nk8UOUKNN5K72lIjN
sdWLbJDrtpjzEuIlxaGCY+OonUHvO/JIk69/wO3FoPE6t0KdLz+YFTeaDPqD+0yh
SZzzoXQ+68mxJTMyTFSKtz27liuC4evw0vHZVkIpKjjgFoTvzEVS5MDCLcDtkPqM
VyDnvPkKBUxtPMZSxP6zszmNabNlP1s5o3DtmNYybR1g4ZmHg9ZrfVYolJFrcYuf
ffWMEGSZ1e8X1+JlTUNjo1gT6OOvhhvT1oNMbCgFGFALrsNCQeln4dw/9nKx4W5d
i+qdbZifbIrues7fGkR9ZnuviLbgviyzlT78tRixoZRZ/a8Pr9liXr4yER9kVP26
WSsg1SjHHYq+G7A3PyoupCdJfDxmb33zwWLJ77qgeLQrbzGeO5FFCTsEvX2EQCA0
jchnoBiuQnrP8b9jW/KVoMhW+NBUkG+0NRf3+ahg3hjDH/l+vIFMIWHGmEwVTGz0
Mq239p438tSh/bjP9EhU7raIhYzMRi5S1/7Ccp3UPTGXWA2Dlsea61JFHKbB3tHC
vq0NNhFQio5UkbGrm/PNZqBy9Bxm4VChYDYZ9+gWS7IwJ8PLys8CGrlFJ5FXwOEC
VxxdyTzQYmDwskqkcPhWxd7/WyNmR/ui6PpiAgTxmQ4nqGBbUiIIzw6DFmBrKCD1
NwbFHteCUww5CMGw6daiw7zA6FYDSoTdN+GfRo2Du+m3AT+4kazYX2BRdFmn7rDD
lNfRnWa+zBVVL6cqkxENZsbtEwucg+sGXWZx0Wo2uBb3rAYc2EPSVz3katYnMN5w
mQOHBeN+dRYMeQ30gs1pVtjWk3lENs4q1FojZ3ndWZmwtN/BrviGx2w+DMZTbOFg
sdfxK6t9miwdQfqCuH1On00K9cTWYdyeNJCLoeU8lxz/gLoqrVUMXqqczeJ+4WoR
g0ceVrY2tO4xukb1m3+XtpJNINPm66FvnaqetZ3GdArPRsLr9Yhfg2yCgTRJPvby
vhwpXqlXlKUCDTOPVzsKSCC6/QrvCfXyRFqFbGj9iHUBOoHYVTEI1cI1Q2EpBm1y
4Du7PjBq8thnReafBxFRipB9aeM822THboO0CKT9YQO5WrBLRQOsMHrKNP9nXpTM
Thgz5vaU5IwKTsZHCF995+yboNA77te5fCHlHauT+Lyu0dNCM2WFwLo9A6zTTMLw
U8gYW7/StsHOxUdE7v9jXoQqDptA+J7Dy1Z4v/nUWh2JxNSXYVRnsbc5XXzG2UMZ
TrIkpvNwJTrvmYyEFRXB9tc7AVkA+29o91T0b6ZAF/5K4Cp+rI3R+CK3j/Rjnhku
X4l3xsxCkrerJ93b4+7aebFO1eYyLCHd/nxRLQfd27bC183XHcBS7GQHGpcQoylK
pC00rUAgiHU83AVtVOcsufkcmnLFSepI7XlY9DbmJl69+MGYGzfczS9QHZU3SC7s
mqitLJsLuXNqxIHdpLf5DLm+6Xyl9T10BWhH3X9vDLuWYO0iP14xresWBYAHBvka
Bk4wNQWvGbIjPywvWCQbYFAMY464W6f0S7DfXgXJu95bVHWYSl9BP4M60PTLIIZI
2n3X9uJK7iFsUL293YDP5kZI3oPT3V3qBmF2+/aMJUGhUlGLfDKhhOKfYVaz8MCj
QYZWhSBaASmnzuvjWSqfpmb6VT82Bc6csZ9Xua17ffjMR03Flhj841sybw1O2l2N
O64K/4/Xw7eo4pwOWxJDhh0iOPynK49FyNTnOjVPaiHfjNkvtYCoXEx5RQnUvQf9
5503eMb+MiHeRJdBqRGn3LGKTJDAVD6v0BzbN/ayWyTRZ5ZnQDQCcAAyMBPE+161
C/SDc7/tGZ4NzZi5oH7CB/hf3y2U6hxGK2IMD2v22ppOpLTMjwtkcPDdjrxhrYa8
wLlfvA2dBYWYCNmJUXiJOIzEft3tmuWtVakY/YodOxTIln9IFlqQw3Fb91fdU+d6
ahzyBIi8YlKRWg3cajURPnORU/W9YRGuLr7lOaGC8qo1Pe1C13Cjt33LG2v0a/+1
zHbYlYClRslnEg1Wnt9MxaQnW09W2AF6jgkN7AqvM5/OE86RmKW0Ilgo+NjQoNIe
+Ob3vkHrYPyLDTBCNUJuKrCsGE/HCVsyg0uuo3t+zl5EvRF4vzyKaAnE+7V1jnMO
evii0VCFM/hCFyOAscvxV323oRaA8OkvrDkach2TAzfZE+kwfzJv1SW87p1lSRRS
BQZQIDQa6IPA0yJejN0RD7qS7ORKBu7dUqh9fWe7qlzR1cjp7NgCQnNlASRPzUZP
vqQhhKI2uA15SAcRau9NcVp6dId/odzx0tSanfDplKm+R7Sd/QrmAV4CUOgiy8wC
TluXL0xtDRJEtVwr6hbHogwPQ/SfWHMZLpx2tRdf0E3V3cH9pXpCWtnvNZ4kC/g+
sPRIl5+/eZMXJjJP0Ms+IjuOdH1AQtEwp4BdjbKwdaU1lNjFgTdAutFtrf1H7vfa
jfQA6bjZk2uJqIBAkXIW/XS85vg2PIA0YbEDA9ttwK149xFKwLVuK+5cPTGZBs2E
soGCA9PrLa4SJyOp4QreHmwqz4L3nZqObF9wjcKr+ZaAiH4mB8v6ohbjm4oGqf+/
xTmGtGyALVIDKzyMDAz7gPiPd6ZP6FHaQZyiPxw09OHTl3+XpVudseU2yrbIdU9p
NSLr3xLsWr5StFm6gLWKVDN+TOcv8wC7FUUkI9/iZTRAifV6oLzdtQ6SrqGxfNm9
jz6eUpqHyo5oBip3FLqKHY0QA4aTJRBdaFXtu2/LdnN0D7sJ5CVnsjjtkmDXFHgr
z0Bf9mSfHv2WgxnIPAPfJHftH5lqzpsCjeR0Gfw+OzpaOFDg6o1ssj6EXGxFKvqx
UF+GLpFIr9x6OezjH2gMx3PyU+mvtm7nzsHtQr3oJKMclfeZztSWHBTDnPfJsxA7
rN/CstQ6Kp/KhOHA/p1EvkgcpNNAWosA1Q6QkI1MKrxTPg82Uw5R+51xb82VitEt
MpUTFuZ/+9xtOs0vdPNATUF1a+/S9MJuJOyB0XXfH57pXE/Bj/sCC0Tk1K/Su8D5
rXHaCe16Fe/pD7y0byB82q5RebkfqV5IGVpScHp4TYG401Npq1StvK0C7e9RIJ7r
yS5ncqkLV6vaVzZkTfiTHHCkcVZO5CplNHMUaTCQBBKTV8mAC4nb6L/Cg658kp4V
Z1bIhDzSBuC6jNfl7O88+8vhQsjWH1L94DyckHLWmh9JRgm28Ygu8KT0NoIpzjrh
6ns2sy0n7XGiNOEsj5nqALj/cZtqJKDE/cH/zHf63NiA4v4b/wpeEZCHV3UdI5eC
kJFbppXqcXaqCpaQwyXGjzl5Z2Rxlqc/N3Go7WuKQdefgku23IQjoCVxUVqO64Yo
R1+nLn3jWTC1a12viwGzQU8J7dDkPrRNFQg4h1NPTzKJIX6naPQVgY3C8LxX/KRI
ZAjZkRIVTdKZYIhVFe8HRNIj0PbYNISXeTWYNBV3QhB3yeqQZ48k6wisEfjQlJPR
0b9aak2ZW1TT1jcBSNi6FamF+Ny0RLzQDdqQDxejcjfl/uoQZ9a/lf7bbySDi8Y1
crVAtrG1IIowG7omk4AitYwfU5cG041eaaR0TcUDZ8Bm0odzs9Xyv+wxk+GIBV7M
HRk32vxSrXF/Uajhwr0cCJ5825sfCVKz0PPWFakRyUgV2PHWfGmFRKQ/qkIVl7i6
B75QzvpgzKWZk5VUQoVrD6Ac87sIH0oSN00wqjhMgOK0d4E6scGOikZZKjKMPqdN
f3OyG8tKlRyPvaPpCmHysvhW31NS+kY4uWbjicj74vH8YnAYcJb6ISSYZlshsfhu
3WiDwRiKSlurfKilGvzctYSW+EuE3v7fwmAVy9n1OM14YSAzvzIQeyaKBxePnOLc
LYD66BTDGYbKF+UYAiHBVniYlUtobi1qTeqf4+Lt9NgaLDtEZX4KJ7n7ts/V/En7
R9CNLSCcV5iNqo7b5TiKbyNVz9pOthC5BwpIM0N0Mft7wBtv0nBist2UbS4SzlUl
nl6wgQKpQLIu5kTYzaYlWLHmT5GeQ8UbyMtWSJdsM1cIwbhZ0sb+qAdUq8snSEi+
66IHVtOc2VM3Q/PQMofY1RBk4s+bm4IvVwCfwqzzwjjPwRb18aR4UHpG8AXLkxp1
SeFvQXf+1rrtgQTbKKwQPq76TTuqF7/AJJlHPGeEbl7LTNAYjWURKmyG3VA17qd4
qIlYMl9a51UsBCr5jxzvPR1oVZ7ObWA80BUSBtNqmGYETbfl1W5aNY0JcA5fg/MH
e0b9atOqD4zblTWSoj0rqQiTBDBl4ZWnB+M/yREcGeGvX4QFael89rZfAlkItbWd
UmrHKNQf3ppDA+M2SX7/iUuGZJ2R6Zoaz03iOpUTFydow9rgXTfLWaYsV6h0Xd1J
z8k2tQqOPeP3oFfadt3ylz+0fxyHSQr/j7F+/SskTWlkTIX7uYZ5cathBrpdSZgs
RtKZUwFVKTK1Ui4/J7iYRZn7RqGO4CK+GhNgvbZz/5dk91XerLZXVgIET9k/JTkS
eT6TNNYhh1fDI0KZtIq2qNJelZo6SPxd2NVWAfDjrSR/od97ldldvWuVvuZYJFwn
heJDGrxljqYg8knjCnrPmaIA4khmMIAR3/wtHrMhj3PNQNaZc8Tm7W5g1RlLzbBB
WstMoGsGoeoV+OJZTZ9AdNFCJrhOSTkYnF8tGGrnsOeUl0LCFhKT1quYemDQIr7B
xwQh4ynEj/nQkojydbzmhSWEMErkRARTP7ZDWQrOK2JOU1oFAn6gThXpmK+OO0tA
FBsIhyYlrRe59RNSbx981jeBURCaR+l7mQ1114SivWPMNN/BhdQyr7rXGMJtkFl6
rB5CreVNiUYHG8FE/xWV5fSPMov5cyEEaSdejx+7DeKOpjjXLqTQpbsf4KCgyFjX
2YboeYUfuYtiwtn+Vdix7cl6XiWOLIJz9ePx5wqKYq5BMzHZoERhL+8qmyfvsj8f
oGXyCbbR5cD5U/6rN1JPp3YRogCpWf6+dCxCN5mPnV5WQs2wXQ55oK2L9p07w5Rv
I3vwrnrK6msEmJJBhxcsBezuWBDqWYf41DnXsfrxUe95dAgTAFqTBkaq0olygP93
RZS2makWwXVgz3aQkrWOW2paf2D5GDpNTZnycaYLiUNQfzDGYhNyETB0m9Sm9FTt
XZBnPFPiyqoO0GTv7hbvBBl+aKKtNEn+gbkgzSXu4mOyzOWV8SifXKFapLM1N+4e
9xpGnTAeIS4iC3vjFXzFv8Bfbv183CcJ4oyfA44+e6IOj3oIRlk8d/3syDwtzlYI
hnXuBIuUqcHGQg7O7EwVwCI7sl1M1Cgb29LolM76kdrScFZXs1CeR7KR/aGuHEhb
TkgBuGFSev7R9fFXgYEfp13QZsZn1EcYjupBeowxkPcsRBmnGeOPXUvzDD8qrNK9
LuRHLbNzJ8cI07DVaeOVxXS1ghNREqr1BF/yaP3yK63oVWqEMXorTMOrf4peL9x3
DPSeS9AfR78NK7Es9e1vCI93csQyQEwa3q4R+zZNRsUtPEGmZMVwND7wpGbdRXhv
HIoWmLC8aDLPBHjb4Z5D9BSUbDukDGOXhHH1oSHyGYWhwK9nMzEa4Lr5egAxELWc
8dmI9rf0Cy7PCj1Rbak/1PqypauiMNzqboLX0bgqMWy5YfKvs13Y/5H+6gcy3mLs
yD4tiSGQorl0AkNaJQ3pcAjVFtGNQHJydHcIS9wa7SKKCOCYmx+zh7biwbF6tJSY
p1TSNMYJWiM8fafSsHu7hDi2laLj5QsFCzkAaIhTGh5CDDw/Lq/cnpte4LbMBTD3
1gxIjlTh1kVTG+jcHC4f1GB+gQo78KnwpAt0SwoxWbiDK1VDz4VIwypqe1mH2ARn
H3Kt4YHhHhiy8mNmsEyF69xtPqvE1HS/kMCy8R8osjhYoxnllWs53jF++nx+G0Tn
FXU6eiBKxOoQ07baFSNOnMkE2PbbW0UGWQrCNweZvOQc9OrOZ3mrvC2n/VOpb242
8dyx0nE7vF/XmUeXZgIvqi8bpMaYDBgRKu/B8/YvEeRXmSo7M2IviduNtoNarn1S
zZr1cNTtTFWsxQccaw6hVStIailJgxqKSVdvuh1kZ1eGIshk1cjhLicm6LXcaveN
lwnum6r5l53nOMapQ55loXAH6LNE+Xh9QMKDj4lY7fmSljInsQJm5axth0R+35WR
rgQBcfwnlQ8nZjpF+U2nHIEv3YjabyGtUrpGfLeo37w+y8neY9ejr6FaJA6+5YpX
mKOviA/qN+vFyUHd0HCUKY8CiTtJpNKew3+ayNY9pvqKSPvcVVpFJOA7F6OqFX34
T0vlaHjT8SDenpC0hgPnUE4cTQF6gOh6ck0dLFxd+RSVl6j9jOjcgNxuYe1M2iep
S2D7p3itkgeryAI9noFdjQpB27mb6Ao0YPwa8KzThMZLwMgZbzrmuTQKawGTIJqE
+fgG58TdZPIqAZwjysOjWqOXLf2lAttLEucB0EMLp1m+0VTE8wo3RKMaRWiZXKjK
paE0G4/VmLOD29SyRtCef0WhCtTxtQRr2FD3kwtPHZPRqgDCbEeU8PpZbbDZsN+h
X5Cm9bqkloV5yYWVZ2vZlNOfnQcEUnDdzQv4uNbFdBHivWsPV0ftcruh39R0J8RJ
ZhCbxtrcAfipL1YTejnZlawqnd857LDjC7Lj72bsE0x1huSFsU6UG5X5AwCqO/ZM
Rdw69oY53a/qXr1AsPqyoZlwfLwalnL/BkLLdsUCieaotbxC6LfAPeatXfnfOF/K
Y7A3Buo9m/2KZiLKxmQTaQQuUJj+1bf/jl1BPXfJPCOOU8weOTIWkijPBtX6vlQy
PdFHBFilKrqHSFNDIMpYqgICcvb2aemxvyEP4dE1/4AF5m6LjYwh6zuXVKTds88S
Pq+1Ec4TTouPB/YlDugR4IOlxBmBwWWwe9TAmqomH8e6oNrQvEnTalcUg5bAbWjX
AMZEUzmN/GTUhF/f9iEXs3KEBifEKn9dyrOhuqVCCGHnlcht2iyDoQIBgzsS8Wax
PKKoc8JcZ7sS+Gkf+Cau/3SsGLrkQinakyw2wJp8d2XtNe1Ncz3mxCYQIDg2bq4P
36y5WVs13eR21BAPAmPJ6pqt5kP+fVchXSPzEZyDclzxwxaDvAsBzbz57p2vK/qQ
cqyFsYQFM2Pwd3ewl5tcS+cdsv3J1ipYwB5pa/O56BiiC3zyodfdn7sDusFf2Bpu
+DIYgu4DMJttfaD0b8tE88Xgf25OsXneVTuoiEn2evi7XEbOLRlF3Ud1wjDLIE1e
g1V2LkerYUVI1vpwTs8CEb7i0J7/8n7yVGXEKqF5i+aMfVUskBtEmaUcvdfzCIMI
/+HWXQvyPc1PLio0r0eb/4S/R1a2A/srlevQYomUdTuseQhyvZ36hYjC/YhwaEfH
08EdqUJ7q0/g8nuPhDqWqmIa/CM9y5YO6Vm7RfM7BSdkRiElggWbwLsq/UwPKRj4
9/yXPJGzCupgpafRP58g9MXr8lcjSxlwEwE8J7nnNg1QDxKIjus3CFfBTo4mHp2e
T6i8d1SBYyETO7tsvkcubU7NPsyOpTziZ8S6f0uBqOSP2SZ7f6DLXohTr1Eo/TAE
Mk7Yph3bGVau6aVtbuonvOrxcOIb1In0BTGlz6Hsib+2wwvxgzBVbfYty5G/z7ho
nOGNVAeiA2AXlfI6hKrw4oHo9HHWU5eorG3pJdT4tSMnbk21OdUw3MVEYNhYmtP4
oqPiZBWnrGueH4E8vqI2u9Zu88hhVWZ/PE2eV3bKLj7BUTRQ4X2aDCjZpHwHqgrG
pu40Wg1vObPvGEUwQcmNkCw47RFue8WBujrBhFGK2rwHez0gWc6jYKjWZfsoZx0T
VUg3/tpNYNfFANlFM63gItL6fKOIP2kuI+sNX0zKRIn/s59OGkt8MS3P2sgKCg4f
/S+E73mI7IRS4JaXrCCdgDqfVLYcPB5s+ia07IdviLO3tjv1J67myPqSuXQ/Eqxw
zmQ6ItTLs1dawimTq2r2IqKoWw5jJH18khKQwtdtkbhXeDbpmLO98vEfJjusWuSN
zBe017hUdfzS3BfSqKXUDJeu6CRvC68b9g7JfiSdwItDR9GUrouF0nXLapeWCg0c
ZzVdSN5vRJLqSSnosk242XyUomR7nBRQgkgHp9mpxNyrvW/jg+GgqD4AI4xYhHB0
tAMB1YX4ZkOt9ZZLNRF2sjcBsPYjoPj6crkB6svKEc+SDM6rpQmgBh8Cpw6O4uc9
+J1nUcQHrjVbYMJKWPBY5/BZRoeak9NzTVXwKi84b33+FK3MO3/BqAkUwYAhW3lw
pKqOUFvFwE89wajCjSd0/XibAhBpoyuRbE451s85ntE3flnMHI4Dt35xnUiCJCjA
aMHr/hX31dVwabLf6r6XLT8dreOCY/RC1Z6cLqbSJrXdsythIL6mdUA5vixSeJP6
PwYEt7nt9jw+fSbtZQAlmYMeJxSzutycOOv9r1jBb1ccDFJB3dBoHs/8bjdif8T9
qHdPAL87YRVOo3zDKkE6eGfJ4XwUnW3mVjmCKltk8171a4b78ITF5wuG2pyMymAF
45RDbDyR0SW5m1vQqkwOh631S3gMh9pq7vVXJCWbEfTscJjZDWFPZ0Q5QbDiTZ3C
pMujnJFKSTpxC1EyprGtdZI7pkmeYSr8T5nSrnZ4CWwS+G1OxCioGuB2pQrQWs0i
GWmKYx/mfzCxajpr23CLS0G6inyWHRgxd73+IewrI3jJQzioVXL6/nMDyQQHB6eU
F3/eLmKjDB0EvBZLbMSkHHSa/PnKlg0yHgoX/ZNNTYvxTgCo8EN5zA7AMDsn72Hm
5amxT3V6jvl0qYFkiBJpG79DqaXb30VqhVwWL0urvzrDL8UapN5xIMFdatEiOD3p
CLyxt0UBxCx2/4zoc59D1RTkA0nyP6PdPagTPL/Zn8fGpbAoYKNDwwQG+dt8V1X1
vwASroePmnAhT3ehPR1YTBHKW9Vfh4M0+guweo2hA1WqMsQkTFCTrT78riYWqn9T
UOpnnnQcdc/fWtiqzsnPdGzD1R2r1RzH6cwBkEq5Pd5qcc2SsrfkBHVtPesuaEjt
UYZmc2vZHRH7sEctsaZ2jJBUfk42QKbLBywGMt2NqjBEZTDaW/5RqgQgmvEcF28t
tGIxLURKA2s1n3AxujtdasG7WCU9aqzRJ+rHUSW26ICwK12U9B5JFnB3IkX7Tir5
5pJ/VrpjwJeltnvU+RPBUqaT2SKFiqUXpNzqu64ao2krXpUvTI23F20na6BntVxE
S03p9trMpfcjq0z2nEDj9bXYjJBlziK8CLOoirK07pM0HcHE4Wpw00qfTAfaoJjT
BRntp5PHE9FVrfZ6YySqyq/hujyspMyry1NPh1R+hJTeORgUOumSwCE57mYDoGbV
r2Gb8N5SW7jEQArI/KJhUP1wL5j1YJ8OT3ShPC8uDT21wWFCJHg2sAeiHismKHYa
TSNhiH6IABcZ2sMlMHek9DwdV7n6ILm0WHUHexRV4EeVZP0f9CwnP8pTQorxKeYr
rQ4D5YGCZpgcM0rxHK5hTvb7x9OivpS6Pm651VLIO2gORjQKUiGuvHtGTcMdDJMw
0k+0QyvoHf6gxQgINGXFfj5GeVSFcBRK+xdVORZb2WIn9hZyFeaGkEVcEABNXt1/
SJRw1k5D7141Ihwmg3VUhQ66Oy/erU+FKnzuhxsLalvvKPwPrZ4Xw9aTpQ1mFGBl
R1aDwijqbvbwIoAxpIgTI0QA2e6jcEFdN8qiCaACx9dO327BbX4BScWbnYSfEKZr
rsFP4e9zfUZMR89XDsurY8w6o53J9x5QW0LmpuvPBj4Mg4CEO2nl0KlcRcBuJ2DG
Z5KuyfyC+VptM5ADnoxc16drnj+KzCz9iKyJF0x9/ucj6vuJDRUJaH4C966IHJKN
3G3cJ6dso77OQ/VQ4ZsP3o96LVttm/OIAAueCfHBz8UPMlbDTBPVUY3/Y9Xpqvow
SVT+cFuNEuK/AI/yR9g+spVFT8sbtA+Lw1XT4OyoMao6Xb4+zUR/UUwotCBTVoGP
iyjf30NdnM+RT3z+7/a5ZXlr6S9FIUpYsRF/pFKu0wlh+Xt2/mBK0jaZ3jApo2PK
oZYmtYzDTrDDYLx+FZ5WyWM+0VY7YxwF6P5gNC+dJg1BxKRNniHDxsdehi31oc2j
cQ7N6DK96Iq3QviOqd1GEHuLWLdBXxWfDh4RKzEiCjOAnAOLHNkLCbU6Qv6/0/iq
VEdwj+aUp/yKFBuEWiJHbv3CN2YXjB4W7yjR8cuIKrVJzVfewYtpJWKrQkILZf5l
B3hAAU0VegjVgYY97nmD74DTWeRmep3HWxFn00q3VSz1HIOGNYQKuxpWKUCrNjwE
YxhFJzN4w0e6pXikXb3JesgQU2TdAHzzQpgr/3uNURYdpcGBtHhKcld14FwAEZdd
6Uiyb8nU59Q4mGa6OrrWmIBxADlXt6+LQDgjTQZKehDsNcd4tERRBX8r6kiZXcnE
WbteU0klpPlBnxB+ZCstCiTyJ4majZHcvd3o4tbDU44Ia3/8zIp6iWS//wyXkQUE
Q4YbNrpeeshCG56I0pdObiPiz+R/rbGxbNYHbrRo1i25NTYoke5TDGlvhvG9JMNp
psXfvECIiIiaxWcoVp7dEUh4JIDO6/Xd8Y4f/IPgs4LrTNp2ZgPaWrAPDZyqB3gQ
x22MYfIjZxUq3d6dBEYVcIEcuaKpSIGNqgb3Am1xiwebVk7HQX2gu+r/cavDIlew
+EG54tnTWOLmTLzsMzxghyDlwUQrt4BfDJZLfgXnc5aotzUxUF+387VeP5YqxPCf
B2uXEQ93ZCWPTHxQzZEiNmdcpewRMB5jkaH/nU6Z1lVCDwhux0iL3RoTCEC4BDJV
+odUJ1c/sv0Npy21y0fLk+XBkAcB+pkgzgM70yTjDqnrCwvZS5Rg39G4P6exH0tx
tfG6Ls4hTAl+ww5W6vWgbvDbJ7cZlkFkD3ha8dM5EtS8Cf+pvJ3eO2KQsFZNAClj
IFCsp8+vp38eN4O9wd99vpwxjtaTsgc6SZZyO1UBJWbXAB7Ozg9R1SDlyvj9xdNn
yWRnW8n6i7jkF9gPx/s4GqkrLi5WDLBWz7kF0d91te419IZWKuM0UyRh7nZOsgTo
D+Nac3BpzyAjMZIg30FAJbMqKzhvOylkM8c8NUHmu+z1qOhDon7rGwxLuVWmkGyx
3cbLH1g0dPou1U+Xt3IJ/cR8aa58X8RUHosBxXgF1oPkefeeRXK0lOT5Wdw5+2fN
O4c35h1QcXycA+AGiWbtcyrb78mDQ8+uXQwyL5cQQkxGv+H/w9uSkf2IgIZFuP3A
b8Jfrs4XXxqe5TUycgKqQ/A/9/Ni/KYSdw8ivjfvEYaykcTuN2Pj/FoCblJI6LSh
rW5PFHUgJTCNxil9cFwVmchpEQXDJEcfyW1Jc3+iCM+KxKCS6R3yXiUg+B0HXsCh
X0rSM/l/IT42dx4cMlEm/ijn8496RTOwfO2beeMBcxJ95lKF0giT+s5gHeMI6pPB
Ptfze6vrvcWbWhT1oZ4NWS/2qI4cUsUe+6jXu4R7uDleOS/l6Pdl9jMKpGRcUkpp
geAV+ISln02tFcBUMQUT0nod6TxNaKqe5WMCS67qn7TQDbTKgda0ewChqFfyfZQs
NIJzsQyGQEVGVAd/6ttwdqNs8TXJtmRSR6J9NEye/E15Ie3ExAQ7xELYs9s5A5XB
1QSpu3QfM3tgLhgJmP7vIzPK7l6aFghnc7LeR03D5ciq75UTqjYosOQDw6aZc/la
IoGthlDkhfZS03MyVaU6C2LYXFj/tYVCiJq4tXEFdU/eSZHgm6gVvbUbCWeM+QcO
VJhRPVA5uiNEXQ1aluhmoJt1DXRUzk80FcGLFEAZpML3/twBw2BSGEYkYPvkCb6A
boW/iLZYNY12igEk79Dcutf8q3PNoHvIu3BOOGxWSCGiJCHFpUJjvmE33Ikpq33c
a66W8fq4wBj1S/2ilIgx7jKOh0Iu6y6RYl80n9mhlgwRKWHzOsiSCSQaeBSlIQTz
JfKbr4Jcrvu6uuDLgdS1DHDyBIRsDMhhHezWMzgnKodA+Nf/8Yd8giIggkC2oADT
p9/Gm0uowBDndrEL4huSEuKNLGz2Uj2jMkmPC8Y4YO8h/AtcyH96OTqVsBu2WZhF
zuPnoLKPiMHvS5pJKzGBygXxVyBGDKAgJ+KXMhCG/8DVfGsLfTh7FlolYIGO/Htr
e2I37gNGfq1yb5D8ifhrWRJF85c8eelOx1YajiWJ/LiQJIZOV8zILWbS9PZxWz+N
RgaVGTGb/ZB/tlQ7TZq9u5bltGpxGhr4IBeGSL2CMHgv4CfaCrX4EsOh4sB1BTFf
8BAeyf3x9HsN4sYLPnBG6hJmcvEOxVTkVYtVpa58b3VfF+2GMdUhgwA4Zst/grM4
gbg4AOeBrD47wWuRJbV+eb1WqU+u8rU9I1qxpni3RXRTngNV5v+s7uormOlSGcIX
7/q4oyQL3jS9c6hI+3PWNvT2TGExYJ9zO6yGBNu0gzKFbT2KJVcHIwI1kVlqazxY
gQXv1bAP0FHtTvi5q7O6PSxbIthaq5fK+7lFTyON/b2U1AT29PMvqq9kwhPtjgiX
QUrLIjaSF1gLiLVWJHDwP9c0sdKE57SURnjWN+rTfx2Lva9JaKc5W2pqMf2gw/mE
xT6VQ1lKdNjqHTNzfgzt/yM2N82u9UnAwveH7X4K9ngmnU8Hr0RBPohm29bYZoAG
J1zTcvupMaVmkYCNzZJnQeGMUw2xVfklgDEgAXbbiUGPfBB9ISJSFYv5IlEuJnrP
ITYGmGH1YJS71pqwVjzjkOrN9vSrLo3fmThdP8ovedjhcDu0KeFRQF/lbgmWslCZ
mDZ8s/PE8pmBX/JvTMYkkBiTxOW1J9f5nq5PwYU+1g0lbUTpSMoOtHexRLY1/8WA
hV/J1PPECpTfOsJGsNOKDweDE2YlEWKAOvHJl1VAaNLVoo4Y4g6pVCc7OuooPinX
Krb6NGt91R8Zh/Edz2M3SrQo7x0QAC05FTL+IqTrJChD+bR7SmCbe/hglQmCvDuk
T0eto1aLEFYOD7Ga3pPUCxYMKZFduToUMk72XhPm4I61/+dIEoIYoLgShbq0VRTB
aD39tltwtGtuntfqmnaz3ibOQIbL4wxjrl/oM7o4WS5PGgCOsfFQCE44bwqE9cNm
2WonKZKJDiC6KXN6QAmMIXy1cAoEw/SkZaC8MiG7o73pUcXyM6zG0akKFcQvmjZO
YF0Mqq18Zak7Gkj9yfwfuxqdEhdEPPRLmnVSY9v40R+hy2mA3FLKLwbJZkMLeOaO
QlOngEbKRsykc+xGJ7gzKBHtEE5oiBfiEUrZ83D8T8weDc0zi6Gv6YPTbQVvb9mM
LGWEHgB6lz7p3mUJ1fxc7IWZH+40vtWaryIcol5hiYtpp7bVXZF557/ADaxpw4OI
qreHO+qGIdXdXEgsTkGd8H+QqpKb08uOZamyhFne0jRHWzDy8tv/3qCjcNGWXpSW
/RbitLLrIqBk3vfZnyAscdqUXfs/jdqWRsjXbsG0xm6lRH62D0XGdU+UvLB/XiJ+
JkiADarMyok9iC4ZKYjFS7zDsaEgl1LMkJdy/pb7jns6Vn+qW6QlIdUDubZ2p/hL
D+hwLO43njKF30UNcHTxL1/UwHYpi4Mk+0x8bHuVew6zLwHgi0Sh/QqmCANQJrfR
GPAwCfMbbt439yY8IQcmUCaENlrRE4icjw6h/qJttVvCpW/vXnga7+a2Yek6yXKT
gt8Tk+wy8g8u6ssHYpBWqFY9Yjz022FlAV9iMK80QUxM0OQcjjtmeHgcwPuSXpBV
8U07MYde2ptZP/9rFvube1H3wqVzrpqOY/lwCYaG8BLVg0PAvgw/iLcfDaJF/twM
uAR6gD8lJjrjEvharysb2io6VQhCAbiziihZbkQWVFGWqQbkicguQg4P7kjE15pu
WMYWEoToSiv2JbGcNseuyDWnnobZ+Z1ZAYYV9FNOWSzRIB9R7QRqFTIxGBEpsuF6
npY8951L9fkEdIye5EBd7OwIZ8XR/m80+dDoApNqJlCzxokbYWq5Xx/KpGv8ku0g
5Ps24pDnr0DYCYAVdWH0JXop37lvJrG/C+9Mj98D51EDbsg1zwbs7d+kJ2WXnJqx
ZR9up0KEFK+8EhozWg7qayfWPi3Alk5lCSdHXAacp5pxyIRJLrkGZxrSKVAh6FaS
IMJjCftoAlaPL2HmlNp58SD2raJ5/S8LEQpszixgxBMCkvWKGC3NXEgRdo6cNijz
zoepLSYiPkVqL2bkyiRPRRjNged00mZPh4Qq5Co/p/gqATHzQ1Zz31uQaQAj1P92
yEgZH7fdfsqxKBeqBFh3IMtL2cQgmHwkpqJz8kfEFiVFR484pjM5Qd+yl1NFcVJ+
zxmer8MAOcPt/AHMKtxJhYx6ooUQEJmeYbqXcGdxJSOsLWsceez0Oa8TNpRYcai5
7NtYVC3t7A66pTKgy+AGM1ED/W7tyZ5vVFCVLHMWvjp8RxMgeM6JeV3ZEClhBrl6
zVwx7i0q61uFQ/F8e+HHGlq3WP5nlxDycpMKrzHqRukI19LIv9ol61pjd208H6Dw
N72z91dPRCeGb0NZQHUCl/a4FMjBeR6Lh1p5ULb/YP5OWwpBfPeTwgclYUqus+rP
olZ/umZ13/fHZx87Qa5SmQyTa7X1zMcZoRZS4kwONJuPh8eWQ0angMH73634qjG8
V+ZcJaHGz8bCc7Ybqm4Op3zVME7pCCxsvVJ+tUvDBYvdKzWticAqJ7S60xlQ+oOG
V51MTdb3/f7BouiTqz6JeF9eTZaqE5fuyBC5oDUSODQkhbnVvlpBlBlhnM3nXwn3
j9mjCQTV4LeLjcbsWGv1VnXFhuoiX0lTMQFlyzSC/gNnwqAh2xzAHYPnsrPHgXn/
HHIOzUdSDIU4fFM7yAbzYRTsERC4kn3hh1vC4B0l62HSBrA52jMguZLnYoP10OwB
4CI9OGxw0IX4XyQd4hVI1zZTLZbHOzu3wOfO6dWX5Bez32kGb0GRuWPHl4avjllj
f8wRZitNxKoOdBkQ9bErxAgnnPH3juPby8fHIgiwn0S1Eoz7xFlYJ9sCRPNOTM1F
Yc5sgfmVQCDMV22w01wUNzkB9BHlTHESU7XPqx4x/KpshlnQ8am0h9NfliN5CpAE
c+ShOKzMAAScJGrrPolbYlcP2vnWt1x6aye2xmBXvnZwJc4Eeun8/3jn8TJOsjC0
AI14DswzU9HM5F3fOiTG1DGmOhnOUqScQD44Kjjc8UDwT9B5P/uoivoBP3eMaIl0
rArVZw+NZdLig0Itz+nQSwdLENyOMrgHCIjDicxvfhojw+dayqeu3N78vHa8ITBI
CRrCaWCiT2AwmhUImhaw89pjO2GDhJ/IxOQP+b/TvUFP23KMndhsfD/InM0LR7W3
18pJC98NE4ph+E90EVbcIYYL3GA1X9NJIYof7VGlFJ8qVu3z09JaN5PEmaxnsbd4
//AIr8tmiLKLdXl+GtZxXB74gkVlJogXA7FMPoE6lA0hZR1W51dQAMBEiuw4nMNk
uAerZMKsWDeVCEdHMQaxV2DykBpTAR93HRQaDwaQXFbCWgdNh3/ZkKmKK29nyw+u
mpNr9esFfAK6g2ORXBaomNNUnUVxWgAAPg6jaQ6fUOXvg0JdLr+cU5XgJF94o67A
bL8rr5yaWl2o4AY/xbhsp22hR5unkx9RVRFhv7dQc9AJSW2kw8GS0GHwrPZihLBs
kIsv+dYPZGuvAbJTUJ0/yj9gVRB1JC3pAJjhmPmUidWEt2NQqfPAny5ApCth53Dm
4XGuul+l1K/RvDaWq0XB1tUlr8b/0VnERoOLfz2qbjPlPU6AoB3nMMbnZl7xCSTJ
aaJoGOEaimKTMcb5iddO09BKj1sHjVcbT7TUh4E0z6lcb/0k+F2fC9lSiQTL1/aT
0cSzIdyLIZ8MTEfZlI6sIgMnXH9wKLxuU2RXdtam9MWSrr4m2zfMyOh32FsSPICI
dfzXab4oyz+ZOsdZxTzAiBvM1nIN/aCjBsSPy3LXjS07yp5YFsEgWB9ZMxCZX+wD
8foAnxwGqpemkXLeTVEegV5uV+YhbgTpRP2Dg/VeCetCQ5a9u7ZeyFmee/VT9bn4
TJeUwDQBJ42Q47zgwu35CGQBR1MShyEKUvVEodnSRY1Eba+ybUfJ+F33fs2LXkWZ
vb3b/NBII3sIq9LX5BUY5XNFW8Jo2uolcUdkJzrBjTafZHA6KltGgfQoo33j1fFj
iU+QqfeSC0/jJu9KRuGefsVnFFMbRvCx5jlNv7xQzACf0182HyRyHemBCIPJ6/Oa
ry5Gt7NjJvRujT0RZ0BRmXoUpjcFS4GabHg1k1G8jOCMCQKC0d2B8t7+eUN0L80n
kIdp5CYytnFmUdydPCyYG4nAvjNMq80gV0Th9mVdShXTgGEp/erbIHoOe9oO88VK
GiBSv5fiw5Zwlyy/mP1JOEGI0fHMeQlKGq60dHHk7eUn62VtdcL8yNGwJHDUxjwJ
2CTPEHH7FH01cFUbBPu7hkeSwD9VzzH5uiMZBl1rwQLOXSCdOT0MZrOtpiWXDpkJ
MfFye/zj64zm63Lv2cqq2bVRMehPhyGfglzi/ZdFe/PQ49o91wBSo/k9BTCcbBw6
+5FCEumQYmrfAMoDjz6ROPyINpG7WR9RlQ4JDqnpkeC0MBSRyQXICZeB9PGWiXxb
3p8tdeaAOoOGx/OfykOIujivj1+gzjG5QyCgPctIumBlapobjrEBYvVVqIf1BHWk
a/smEepcNzkJ3Lkxld9O34clrcQdg1R2PHEUtzZkyOII1bHGcLSP55NbHH3oupll
1llpWg2sg45V9vrCE2+k2daPMuiLC2ZovTLPVJHL44RhqsAQlVKnI0FAIaATTOhp
GOczypbdlS3u55SuQRDvWL7ujwP7hFO/TC3SBuDmBOp/YwM1qig6mh3oVCVCN5w/
QDRSc9mJ/S9IiQ6kAsJpyeqesZRm5ghE6yvCIzYcAVbcnlPUQeyoK/vGx58MlNr7
zwrzjy8rGtXPtokZIydM33DyM4SEFYMbfSHNktEQp3UgSw1u5QPRu+ysfQPN292i
s6dArjw73i0JmMXPeGJh4sa5w3feWFTD0aJ1QY55O5Nmfwbu//NUuD53V4qNQYvY
lNhza3ksShdISkAEeoZDtiSC1BT2x7yQf3g8XqsRxNZyWjeZtb+Hhf+gy1L4IpWF
nilG5Ko33c0Z+vtGNNOmfPBRYV6i14dMv67pATh2skkW38eWFKGydPiABEgpAcaZ
RscfA0jtkmfEZzDMi6paEzd14fto5UJrbfAUZsjyA99KZkel/O6gM6A6/NkbWC64
nsimjzYfsohhsFA4cZF4qjHjcdtYWDFLowNhjvUtV+pf41ml80C4vvV50f6ADISb
9BLJNTMJfT1Vvv3WYl6GlS79KsDOC2Qlriuy+ndfuhVAlpO7/kJGNifoH9d5KbVF
T70CvBpojTjcHHzaSlecAlnB/N6iS/2LlVYsX5nApTaSwB6E+VC8jWWItoqFzcDc
uoy6apW86lKILIktIWb6KLJ6SERODRaj4Kjrsg57VunKC1ftBI8sO2q1HLoe72Tz
96iOtRoeF9SGuf59BIDL09ZVhqegUGvp2nRwMcBe1HbiyJk4PMoSVCEUJ/jW6Crk
b/wurAQZd8OJXMgdQVHtmJ/zaDwMMr1EWeHJUWNut4NFWi8RmlkZfi3Z2cZTWkFc
cUkJ+Do2eZyt2jsMebNo/KMNbBJAUNiAbaX6Ey8MOqX13iNgIGLDAuMYZZoE/5WA
SBPbI0Dc46PQfg2tX90A6AMFC6NG6vsn17t7btRy1NbQd8FV/7rZPI2fTgbS8vvm
jURAP0F5lY/UwUlfHJtAtsE7fBNcuhNOJEsX2LyLAillUEC4oswVxjlxueAHdgzI
0lEUgpcg1KMbzj3k89HbAdZTeBni/YMxbIR2DaVFb7AH6aFQcm4YZanMEQEvLL4a
9h0bZMiTyQorVE7bgLoMSw9w9fJYpqDp3zkq3QiGXiLzUKICqbi1Rx8U+CRJ04aM
Eoa5xq2tceU2OP3lUPQeU9li8J6gSAfW3l21T8c/XVSd1US+F3fLxeXpxo6K/V3W
fTz8GEIoOOZADMxCmslNWC20hW8mCA5LH4Zv33xgPeeHmwniDujbKoGb7gzwsAmN
W7VZpvVjqbonzMzFJEwTEr/OzxCsREeG4AIGV4+/KglAa/1wvVCiyBGZMOct7Pnw
gxpWln5KKTPFDA1UyKIZbUtfVcVJooYxvtO9UxM+IGjbZ4BmbceeogvnbwDcFkgQ
cV+ZZMclF6GwOQp+R3jWOR5GwReqUGrrsnubTohc07U03Groq9axbq0KgMZWDC3J
w51NeepR9J8aZ+2b4CZSfCiRssJ8ia2F4UDM7IBN8GIaLBVcurNkxwdjqaanrAOV
j0jx31myUkF7Qnlf6WHRzNFCdE9+fFeug3FWOm+kgFvmCQYM44Z0EA8FO7jfJOSj
2znvRcIIXfeqXME2TZYZmrGkiJHiQIBT3K1j521/o0T6bCxF/YiEEdRB9wrTP5FR
7goLwEY++1AW11escAFl5qaeVNivqmZDqvhuNHQgZuV5W2690pL1iJ9xhoaeov/V
YS5r0M4iy6FUu8YwfsTrFf9+k0k9m/azMQWUxmNfEG7fLP1xPBrPcXG0jtUHLcRL
0WwDJqF1ygmQ4130DgwWEFbXHIwXesU+t21CilaVEOI6Zp3Jd6PBmg5r1y4RZj1L
S9yNVgJBrTGbbtjt5BUaaVdTvXa0Hhxo/e7Jbq3AuOn+NxI2MIcyG59YXSDzB15C
z4rD9YK1zaYjRLrzJaLYsfyreumOO+8Q1cCJkAmlnYNUKxa51ZRl5Rp49K/Dl6z1
+BUsLJpn+w/ttJx5wXQvgjD57884PWhxBjMDrbjB7c6coDqD6IOmPpRmAVE/jlkP
UAJwng5NHtl8egTpGwMueIZra7nXQQEgYWWCHtT6TlaajSFpD9bprTLsCMI/CT2C
ibMqm/JONcwrzf48T26o0TcEyqIGs1gpF3OXjW6smt1J7hexbZyAaPMvw+uv86Ua
yrcvFth0JpDn5bF2zAYKzFuNUu2Fq/OIgXyhfN83Yp2P7e3yTW7vXeK9rcnjTJ0N
XwcQ2P35QakIC/gf3aNNjCWgeqPza5veKQEEGMZ0iRN96UWAhZIU/I0P+4UtEpNI
xbG4C2xkmGDa0g7M/NhnWzM5fL+Hr5aLdjxhphm/HoCnj08iZATHSeKAjj2knq3o
DgBDKVmgrsNr8/X/PDMtvp1DSz3mD3V2+anewHTSSN+Ov/HBDrKZ+ppE3qFc9zZL
dvfNVqBbjjp7kneFqiF0VRhTbT6DuOuEOZVcbn1PiC5wC+2nPqWjL2FkCQkAURL9
IjiCh+hIMqfeSDBj/BHfNqKYgwtlx+cdt7rCKkKWumaNkG66MADRETIdJusJqgJd
e/xD6X3kbhb/r9UYuXa50hG+x3P7wbJjfmceAeWJ83taXBf+jQQnu/Q/xNnqDSXq
Chad+EypaN5GYwtvUZk46cRGxm6Jmq1DmTbJEMfGCPLNcOwLDYvJlYT0IK0MXupS
qvs8xFmChaOehwzeZwjXLTUBfKWLxxtHn5RJHwGRni7aaXlvqv8revy0n3V1MPCZ
8S8PVCuxX1mYjmmp2RCdxwTm+fYJG+7HZ2UqmndlaLKavN2ecZh2zSi8ohRu+4a+
aiQ31epY5hWiN2q8jXphVhjYQC5eChdQ3gNOCQwM+ZoQ33x3gG03GRK8PmnrrODO
LOw2J0EvNPGTWimnvhWeiTMAok1aIAGGVYH8a7vmzy6unz+CYgglhvluNgsdtb1B
fwwzTX7YFdNd2Ajpl3kBQr1PMCrE7pkL23qma13fKXJeGa/sECK1n2wjuZwOZidH
nkY0wwWxg5WCkuLoa1uiNNACvGOSGpGSWOzBwlI4gXrlte60qXUs3C24KMW1Gpk1
ku7i/MVQEwG4DlHsjCGq2NH5VJEsEJOGuxuvtyTzziFSIKD3t7agMwI3tC/JuVPt
1x4c7qLiEQ5iY5a/slT3z4z6vnKDihsDVcDOPc3udZc/DjOMadiFn+oYjB3NNlNL
esY/cvr8/xbSUOswhxyZvQ4D2qjrlOqkhxpVFrvm9tEH/VjARiSEzuQemjzMGsv/
1uaiWXl6CVgk9+lOI8YdziP+RJeaIPTtRmVVXE57F8BCDYT38PFHoiWLLBABsHLf
Vjn9VRBTw6NMAEnSDp+JRPm14O3p5ns9zE48NvCSA4+z9GeNoIpv3HW9l8B4kw7v
9xx1W9colEIDgoC7nJcGKyjJ4d7nBWY3dChhMxh+uZD18Fk3eRNJvlfIcM3aWPsr
pAu67PWHDGBRygd7/YkEYI8a0J+WXBG8xTO87caTARCeDTzCBEnN5qXcIDO77yFd
+iXl/2rE8GgVd5VW/U8/aVbQKw4qSJCK2j7GWWLvcWJ2Iwi8uEU1xtHmmDUhFOs0
WDeDmK6H63YvR+1hG9qruXHsOvhf9QX4T9TL3RMNjwJnbxKHZnOvc1PS/woLOQY3
YCiy7uLMCB7mncelS8g6Dewi14Co0e80dzjiMqvlO2xY3N9Pb/jBhn58VyUm6IZE
V8wlVkXeMOJN/tDTcKFdKpSi+eiW3wDSrXuRgSM3plRqkvRZDdm4QMfluDmOKCJC
1MXvbNNZIMjrFvwRmbk+yuYYrWaMs39LBI5sZESgddZ1yQK53NM9hk3KZPqzTaG5
oBcnBW3SkWtUFt3z11tGHV0ET2e1R/lGoI3+QGBUWnnvIHYEASfKrk7dCWu0DLkI
js3+ercOpAfOp0F7dH+FefxXfKWCJAdTuQgzc+JcXfwdb02Ljq1z2fjhAuaVHffk
XPJfL7cdHzyEoMJAWNrAovbz/fnJ/mJsDBBi8Fx14XvbeFGAWFvg3eETQQllOPU1
FbQOtEGivuWAQlnqXdebur5pZiXj7YHeNBnzP2wPhfbJ8bDdk5+rVZFVRibSn7PL
5bs9I+ucneWyczikorPtE+LMyTNTJQJU093Tqe/EmZsH5kXDJAD3fM2jV8Ii6uIK
oLhuSUVCZV+MQnSdgTmw3EjwO+vNtOSNITBp7QWtqMYRWCeaL/Vap+W4CngkT7h1
StKZ+8adt2tAsmno7zw64CczDJjWKx0uzuoM5dMppKYkQY1GIEmmk2f9YONKRaXn
aAS/35bFUmA5jMJnERo6M8yv+WUvAiAZWD5qDvJr9pXdCLierIEDq5zmGNq3bfpu
Ybo4T7NDHmTYa7B2paGM0gFUK5KcX4EJbao2KxUBejFuRgXMDtmgXMDQK5vhHFYA
EU6QcGbT5oZpUmsaYQ4vpARcneNTzV1SbPd0VDOiV/WE8JlXEnrMjtnXzSFIw33t
2phrzu9vOjgCXRKXQ7ngCgbK6oHd/Sk01wvKOrXlGqcJXtY7Av8bw1eckJpqyYJ+
ICgW/eu+cp2EvSBwc2B44WB+FEPG/RdI/NthzgAdo/idEcds3idNzGuos7z24gmZ
yfGL/FXrDWptLKw5RB1wnbNf3CBrFeeH+QAmACsYCnCzdzb3rEMs00OKCQ0Cg670
S3c3R4c74Jwo81M2Al/oHXob84VV1Zai4kpp4WjhULQyfTu4rufIbITNQfGms8bX
GmIOa+8ygM/v9Qzvul6Hnmdb748kuEytunO4BIP8NTOPpdTDFUYu0FweK28xTJlr
vuLk4dU3niZkUNS0UcyTwzG36kOcHpz2lHVqv/CS861HCvpg8ms/vzvx3LmI121R
8NlbE7AmLCevvCDfYG5kmogSQgqfuAH9J+vRYFbbWSbeaNDWT9js5eu6nSx3q7zn
EBKOZgTejnkwsS4KT14NcBrSPMTZ1kFCNvWcRD/+QZGS+Bu6mqZtJ7I2EUa3flPs
8MQd19xklw4P6nO2MxYNUUFhcynEXksRkX/MHq+BAF0mrtfmxjPUbAGQX9OWcM68
+Au5kq9Edp3kS5aa915J5COmQEQ5hvW3Dd1ag2An8SWFUqj4d+x4YtnoHEgu+KG0
zVCt6YjkCj5rDVrhIHDm9EOrotfY5kgqmIB2+jYsgVXx1IjyCdxNFCpqI1KmjXd3
Ulnjk/pSTU+wq9+GrEi1oCOvz6ulxW4d2dwdIMWySStwms6MfI/GiBeKzZ+FEFIf
F27ppgEoXrefEBhPodGO4MeJLxSsVjulgsdtD/cQ6IEkthld2vzxZyTtImRgFRuk
CnTKEV9LeMu22sHHzd6EPnFrUthOc+ovNthV0wQ1ECYRprbMqiZGB72PW3G9Z645
lAgzhhuNBaCIadpmyF06EeVLsEXgI7Rm/oRGmetftn1sWZWk/d6LnqFWHFKFU+VB
7jGJAnxsZjU/jOSOH8D7J9ZCG01NJ0cqS4hQTjirm8IoXolTr3hq7CSvgqmee+eU
jwNpee+jIVeU6bOF0WnKF1QZ52BV8JaONDI3hICKcc6wOI5SDRHMlS5OMisxWgeX
Ne5uoClKvJRVOMQphuSNCg5i96sKMnDqWqxv8vyUfkJo5zukB14srHuXmD8bP1E2
vOaEblsjs3ZImADJN+mSt//xlTxQR6J2Aj6sU6K6xhKkfh29ihrS5xlydOoXk9nW
hi2dSI72LMnszAASrITzPMp2ybdT5pESVxRcQJVxXyFdvkAZcBqOI2xWmRcSfzqT
CncC7kpwmdezQh8Qfl80uzWHrk1MtE9aDuNdUe6UW8TV5DpZKZs2bz1eEy43V6Xf
fE0EumjZgAdME9G+19pLu37MftVMzEti5xKbbBCPpNXrhQ/RX62vCdQhEV5x8W0M
qIYNhBZcXXTY7bwFOjjZ4ANYzjObWqSuX1L6vcV0CV9+YoeomQeUleeS1+kcUCDF
lK418iBl7gBwH15Sr5DuSbaeqmZoPids4C0uzawPS4aAhNjI5sDWLriaux00YhtU
m+JmW362HQNOeCDBN9woJ8fhc14HBBBWAvULMOcmuODfnE068YZwIyezsag4vPk9
jhWpHyAGTIaVnGZ6jEldnrVKmlvXKgiafOg+UckxTx9NolnAo7C6IISzkYwany55
Mbu5NoM1gH58Le3ssjYw88OGag/n44S1kCo9MxIdLTmBlC1N7Dq4H/5Q4pHhGfKt
W7wPHzqfzKiFBMINkTCr7WyX8zK8WeMzPXvSpNE6+zqb6zTzfB7dpFDt3Q5aNWH8
TRsmW+nfZCxwXqRYSCt1wGTooKFNHHrbdV+Z+Jx6KTJEJhZlCvJ2vL6K/k0ti0Dl
E2TR2IniBrboD5cgzHzpZC6NAu9gpVRO4dWBey7crCa3AEWWq4LNSzsmw+ISiP4E
kgmY+fJqm/x2hiIb30Yyr6anXRqJiDEH2tVnPCNNRcF/xWIT2OqLThCn6yn8ZNA7
x1E6v3BO3QZfHbiE8iq+cdp056ZDuOTbu3AvI9wGGXOgsiDtz06Coz+LzMbl70kZ
hLLgyMnhJ9IuKG+DrczpFCtGXmy2kNzy/SxLWxZ2Ds4hOeNiIMV3rHr4otSBAPow
qY5LOHPxzwf9JOYGiQcdUDWYo9RcFe6BCXUjdXx0B6o5KIKa1L8tRT7H39hIijFp
DKxBwtATQiSSpLh7pTM2eLqdUXmKs9rJeVnXlCFQfkY705vnkVRrz/01nt5fZC7U
7wq0FnzK29BacTr8VE8zQyb1liIMgoMkwaNNeIeLbQjgVwJZ2KCGRG7kuJRVHdfX
F1tNZzecjRGXfCqa71OJJE5v6oFxHaRUXSI7vtqHiqyBwKj9aMNw+OEiE5+Os/DD
aHrmnThYzie9t+xeiUUfDXWupxW9YYykjU/A0QKVO5EvnmMMspfuSXjDUp4mfKeR
4aLzTGSj9Ugkhu3N7c8d5PB5Ypm1n98xC/4lTCiuXkcS+zAb4s67zs2UyubjfawS
JoXVRByijqqrUb/v/1ZBtn7JAlV30Dcf68BXUs9wYRMLMsTRVIHSMduezd+dqJOY
vIoIpIHr8+xLjCR69xYSGb3lLQoFkNgnYLi6Z3FJ06h4KoHCgV8U7ya73/yXgPaY
mpOn5N9SfQyozLqAM9xgm79pu6z9ybtj1PcUNCtLbVf7inyCiKJOeuGkTtlIVvsE
9iXr+OyWTYjIUJT9ZVgVz7Y3zzRp8+InWzFoLUJgjMckTmpxhe+DuwYpXPYDvBDZ
rUgZdihb/YS2OSDrFpWaiSu67DV+qbISvtX67lIOElmopKqfHN4dqevIexjJB4k/
cNjk38mNakgT2hTJO8aedHW7rNesjQ71MktCc5w6is+ALThcvJNIffMnoAF/w9my
kaggLGakZctG5xjaAbHU02TZmiQU+nr9U/riZsXy2oPxP5cTB24Ws2TM6qrpOyyo
F9AiCb5BOkD8xa+QbmwY2at0F/6xq7jJDEDm9LcEHL6E85GXNaX3KX8z43XTEHyk
TG60Q+iFDLwlOT4VTCxpRhZmgolmqHOkRxSzi5TbTLryw1AVvf7o/qcgE5sTdepj
eug1bXhuDDRiSeWkrFcwwfAGdu+97qygyX+P31+Wjmp/UVhwsA02GqEJL7JSgnpG
ru8aKLWon+utrEL4OP/iTY0CRxS7T5ffVQ9Q6M2xR8s/rOADYDq8jgWmPhtF0PdM
RPwpBjv9VlGgwYYFpwwywcPwKY/TMdlcpQyqXvwqM+OFYtQExz6bvW2lUWhROSmT
pH+71v7Kdihndv5U5mHt3SGH7Ftm78AVVZgSxfJ7Ns+5VpQ5ZdpAi5AN8PjdA7FA
AhrvjACLwCOtKNmi80GKfe8292I9MMvLKm57QVDvzn2oGxkKHub1DCvzxZVEiNBO
mB2siw8rR9Zu5waID7yNXPO2knEORc0RCz2z9Gi2Q852ORy8qXmLTLGyZmxTN44i
aTUe6fLGso+6iHXZVhfNMZ93ejg0Wn/01CJblOwcDOquumAbKsvC2NDllUpo+Xw0
zSC281Ttqv8BPAYOBjDaLJrF03ygH8SO110FO3XoCI0OXj+S1Ey1hyZN4p7d2Ys+
mFthEzs2HwiPqYS5/KvMBk81gPdoTJ5qlNGErh/f6WfGKrYHhingi1wKYkQEAmCs
S8SjW356tc9ezNUkUp9BlB4Cb62k/w3/wYWgXQQvrM8jVAlgSBwF+qaDuxaZzl2+
Jow76g8c5lDOCY9FxMQuQHyPvoMbZ+VA4X+0Ia6seW8/Rk12KUkm3HPnK+/hy/0X
7JjC4VTR1r+W0Z7xU5U1AvZicTD9rennXMIZAHjadEitQUyAmStwZG4lX3VAJYfO
Kvf5I6ftD3MvxOcfNp/B3SKkqDJ/vSW5Av91hFB69gejIAY44Xa2EZea8oeH9Bvw
h3M0l8P/dMjMC/wD2DBDnls2EWgTRXZcHgBVrwXI0fW91cFOiu5+iMRp5YuiUDH1
vsU62CJ9RWNrJedljSTPkrg5lQs4Fd6kZfFKsCLp4TOSYmFjlFYUUQG65cMKozCh
HdAi98g3hmttltdVtgr29mu5qpGj2w0D0fPr9F1L6XsRYw5szHZK/otr32bLQ024
3b0q4pHpdpfI90BLzL8U8jRNjp5SXRxrT4kmskDSXOQF3HWlS6LU32Jj+eOHLYQr
qN6E6hBDWnl2YLxdCGYpFfOwLha0xI5HtS9WPSR7li6LO9fZc3trFbn2polA+mbT
AfO063rlHZqXosT2Om67q4gZ8hr8zz9GZ4jYvwcqQKKZK/gJ05lN/2BzsSJ8NFKK
N0UKe48tzdrVzNvWgTCiQLpyt6II8FiezkXW5iB9+Ymo+TQaCPbe1w4kNnRM8VKd
d4nXoGU+CRgcIfWGMkt3+FxcqK86LcR8pp8VWNppGsMyUOPjG6gpsIOHeMr3qKLi
m+ClVOAlSqaq8Zz93Jq0q2uDrDVdNyolnWbvpwrH/glBu4sw+dfpmjtx0+WQvmfY
xhO1p3PoebXy84eacwWSb2Y6zbnao6/7835Ne3Jdf1/mMeYr9187wQRRKlunGeE8
ykpDD2hnFpRF73d1gVHne+FuXZZv3wYiy68o3B+Lv5lL2YTEWby4gsImC34mFUdq
ZDgZXGBKw3sfti3rFHOb+0Zz6YK9s+FcA9RV8JAPSclL9hKZ3DJo597+1jLIMOUr
N3V/H4W++T8opK2t4vVXiY6Fn/ive08meJV9l8NEXiKcYXfap+mRnUaMfQf/h3B0
8zfu4dy3aOlsVwpZke9j0MIX8KXGgQJWhozQ5uEElrr7ffTjOfF9g4csytSw5XJe
V62qAZ+ayS0P0rP5qi+mmEhGXKS1MDsYC2wqxYbJtJVMR3ohF4RyfNb6kg+k5lpf
L955wYzLORsZA9c639XkiPcLRTNTk60yIAY7RjatCQJUojivTPNUO25/DG2zEz+q
zYOrDfZ0QohC/PL3fCZoFDfPdaKcF3/XVqepMepGWvlk8+qIIg7Y9Bp35AJarcEf
qzu5L6ij30CP/HXkpOYAN51Nm1kMhdZ6FfoTLTjk4jl2E9lA74Gwx66kjKTEc1xz
iig3B9mpdVjuxPxzSL1iltgdft/m3ru0CHPh8MJim9DXnMgOeag/PQrmzfmfFFDM
37Os7dIUQrbSoS2bmMbL7794Qo6SXc3JgYjhrwDHbIvaMF36J4MgvPDYrgeZfXJs
3GI69GtOWOWTiQfw2tzF7DWdCox/pehBBcWq0vcYjd69kHQ8mVG/l0UWh8DsgM2b
FT2kJPPr4W0/+nt3X1MdKUbHPQZv+BMaEw/eZJ4A3W2R0LV4Bdwznoju/hahRoQT
Ib7gpjOfJo6OsEsbTFgWFIXxKlnCKm7b6bqhD9FdjO/NPkmGaqZJf+Te+o5wBErF
2yqaGcGbE+VFBywemgA+gYh2ZDWfknIhXbnJ5a3nssE5ewGMLDgaqU5WInxePhWH
baxE22AhZf8TKSElMhVFW/IBsxC9QhazRD4blxhGLv/L9khOLFHBSxSpgobGbQnn
4+E4yDR7vQJ2PLOswR+uApaIoTuQDdpvPpapGTCK7PCVJ9IZiDRzPpfyz4IJW4jD
LtvqGr/3etRXAJj3pk5ifhnv07sLGI8F74TFNEyST6GydZoUi+0Gt///AZvtM+kl
3mtxn7Pgh8XDcWuSOiyIXypk/s4uzMFxN1FD0EEmCqADMOWAJMDLt/PKn7tEqqAt
B8AV3jo+7YOBvWxxZzKBto20tzx5Ivhq5gze4BpVf2x/Tma1mDti/u4YvBxnfyBC
QLdzR9CpuJKUxeC+QczG/PmEGKdB2nnrzL3PwkxI4gwzheEoGHkElcAeQWRWOMW+
jcOLTPyBYMqTgPWOX4Du9vtlKF6Kx3NMYB/PhMCQXG4hDfvZ3tU9VV/EfTiAxhFq
mEfbYVvt+IMO4xRyIwINDQXgp9S7JotQXR0qy8GnvGh+PJwLhdOcg8QmxgtuZibI
/hU/RfrxAGG5lQUVLAyW1qxTfjMD4tLY6J+8VdT82dGyqxGhPAYbNsOet0MVBY7q
aBnpUIRYc/ixOrS+Gf1w6ZFSmQIoTnfNYQqsyBpQ2g/y+W3V2D/tm+nYU5JVS+B6
wi5oLm4Dmxh2O3uggbbjLrDivuTcXJ9VABjzbPdMhuri0tr1oGaO1arG7J946TTx
T0UQfMF0gxJJDya+9R/rNMeZosCxO0XaSmWNj3WccZcbytSswTI2sey292y0L4C0
ll/NhbjcCQc8Xoud0jqlu4jwzhkCVc9SeEBTTMpCbdA9XK7EyVokh7O6tLk86buD
4UbsVhOPPFJg85CKIspYzY1obxKHPXwJ5bN3zpkFuvgUo5l94Vc8V1x+8RfgQzcj
ics4dXDFB25rGbiFTi9KJi03gTwMsk95L13SQiEZcJoy64w6T0MUozNH8e4ImtRd
6+2YrmPbAkIRRuLOk8FZauXDnjfSOLx/ZkCfPMyyFchU0usAx0h1I5xWR09JSkAs
l0QvxEFlMnQIt/vuCaK7w2COUJLkFxM6qCi2/91zQRACOS77h3rqQYjsKvAoPMA3
N2eOD/Hep/4XjJeFCVf5FTY8yOwo/3IEZor76iFu7cN0wiQ5yUgfnGwrs6FtM+KR
Vbb4TAekCY5f0HMg6hysNAClX+lDAEwEOM6yzOB+e5yH6WdNrYzA1kasF1l3VES0
dHi04ZFw8lIQ3VbOjXkrU/AYfxy426lnmUKDfPWx5LJZRPOm4vkCCVfpBS0RZa6d
u6qQaRK5mBvuq8DJtiPMwU+ylF/R5NFVDkvHO08lQ017EQIsplzjT3jifrzcv55I
cCCr02qk63PWTkGFzcyJGXW0FXzA/Tx9BDLcdGFh0c9KwpMA+Vc/16Qt+NxBjq0f
Q/qnxZ0eaFOimtzNp5b2VGnbxnMf/OFB70IPy3uWf/+3MH2oU28VSamEXlBCw6cM
/h4Fe6CBJReTLzet/8kvEz82DHuHMebRDpyohTC79faWzw+ZxjDB23kX8emCZ6b/
PLTpQnJM+eLT42/pna2waKu4KdGxvDTy2oofvGmkyjGO5K3ivpPg15F3RD5D5mCs
XCoTjKWUZ9pJTXqNrNqIPU9LV6PJkGrMjHY33Rg43VI/Zfw+B+CDS80KcA0y7Ur+
RID51nEePybDSoeFldm7pK6k90/f+h49Wd8k0uLAHIjchYNhvzAx8xbV8hp+IaK5
CvI/UuFSMUjLC0E6OM/VtH9Y+oHTvgnQuh5ZrAew+zzl45j+D0C5AHASKMTWZpn2
2z8EbcESy7r3fitvjofvMeax98597S8PEzNurGBIex20WQVTGjXUM0QfjI/29XcJ
UDUUfqSChCjyShmTY6zr3OSOKwSN/AjvKKIee3Xb0I60iBRrNGRRnjh+sS9URvDV
UerEn33h7Hjf8t4p18+fsaZ+UP/ob3qOzQsXdd1LAq/71aPAWgmETwkpVMD4Xvw0
oK/LmSQUr6Oz+YsY7oRYYLfgV+Xmz3u6LmejVKkxHJLccKPqN/22M3GvqOFV533P
HZGNNrmLLuHZxm+Srd+CyGUMWkz6wM4qYZNeKLmiA3hiuM9yc1Q+cNqAVkogq9dZ
bnRwyKbPOhl4kYyE4UB1UvvdUd9U4RkGJox27vzQ9+BKQ5cTWQ7fAKP9dJfDKgJM
DtyrZ0qujjRZ1seCo31M7JcLJBk2CPFlLDNv6CPw1VJLY3beRyG0Gi8a6bUKgw4q
9/DHir1Bvg1ZPq6TiIZ82khU8yu5dLGu3F6l8NqjO6D+i6CRBNZvUHD6yTT5oei5
exSAc4Htz9rBplYsHqWGjfY0P0mZi68yXOiSI9Wk+Yjm2zmqQ/714/eq1kUAEy+6
DfmYT3ZvZRHA7v+c3n1TISbMYaiW6OOBKj1ley5rZGJp8ze/zrDce0zOsmWP6FxL
R4bLbDfM8tiLrtbLZlZSP9ZA45ah0L1umhaYmJDdjuIXu1o6Rcx0hA1+iPUVolgP
1RPvKu0i7JUyaajwI5I4zw93sUeX7Ox4xpfvvzfDB2Qg6pMYFIi1kjxLesPMJ299
lGA8EXRtygHG7OJIy7dZMXdv8pN+YVVv1K+BfGDP3+YC+tWQlLttRyBj5CiG/Ucf
OIJEyEnDvY/3ikmE1e14O7an72S17iZnUh8EBhnR5oYTsv+j3r+CsclTdJPr49KU
TsyyEv8tsPn3qcVrBF3sn0bpGuaMH1NC1ytDXHctRhlodsQC8FqYeB4zPJCqbrR+
WMmLXzN5hzhsF2LoCgGeo0W5ZHxGkvbMgQ4oNJlp5RGB071ub70KnvpGPHJGPPZV
JalCYoHFBBF1hOs4xizoyDrj53WbEflK/u9GKFjSqTqNtvH3XPQ747tBZ8idjmQq
gPWEr+TeEnfWvOaY0jeUxpzghPKVSGwB76DloFLpyS1uY0Zf/LRUlM5U5HPGS7EV
alRnUZTzDgNtL8cLT3+DnOET+1mQhbkQi9By9q5VbB4WO1odxFmVffRCzgjmbm+j
gj0v+J4VlxQRTgW5jJIF1BwiIaYTBZcSZe6E9CqotpqkT0iwuHeln/S4Dmrj+yCD
9umbPJjODFa3dlI9Z6B86FZTZ2FQNOITqETM+cJaqjuz+VWyxTczRTxp9e+oK+nF
5M25U7bt32Y8PhqaO4D0oBl0QZtjioBbfzcQhGtvUgj7DHAOVADiitf8p23UJiVo
Jz1ybArcZ2qYXR5gGjNITXV9OxtllOPu8ydc5+0jgkfMdHgdDa7FVMjDUQXvUSKV
2a/XYed6MA/RxR5x5siPh+bW8cdZO+lgf2DbE1QN73AbMMMWOO3t41a36Zuz1tNO
nAZXjt5hamhti84QwDogC34/0jyJByHU6oQCU7Nu34tliUUBStS5hwMLy6E13aoP
vIAnNvtratLYd/kuFhYU8dV3FxGStPvV44av9w+mjMkWHO+5sMX6FEiBiSupaLte
CwIrcXeVEU58JmvP11R6cBA3nHKJMweLwbaJWzBKFcUM95EXDbU/36Z0cisFjvci
b3o2oznNcn1I1xnnm5374uFqjrGRnhA/V9ph3lKBminJgvQHOSI1wAYPCdywzQFn
lhicGEelccPujb6tnRv2g74qhRwU1bZYX3RNYrxezjNtXc5uMsFBmL3nShxWImj8
k+OjqvYmD3zCSrEtaf2IfY0NBsG0aJeJEv2xoPFHik7AsS/9kOQYrqzfy8KzntS6
G8UsDEro2vdyMxyAm/Pcjv9OZrVUhUwu0DeK2QeylwNCg6tAfswaYwhSykMzZ1fd
OmWTN+V/8lzse+JDWJQtLwnjzqlLYk12gpwJqgctSZc+N/k9BbNRR0GpHtvdARIb
S9AWjsINE9ujRlSsTITTGsP2qLhw8oGUkcoSxIim3HwpIB80LDjSlnCNtABVS8an
bgPoQpDn//uIXBdtCyDOR9izfVhMKqxtL92RMVgAwPNf/SjguHxdkdyKCBGJgVt/
wL/hE+SPp39IH3dqs+yl5ILnPkzzNsm0ANeXYrToQ3zWytp6JngzA+Q2trYfns5X
bXT0T6KmFGbpnbDSMPg/fwjTU410femFZ7GdYgz5fc9Lhmc/f/Sw+9QadQsbrmvD
zhCMgJg11mmYAoNnW1VuDuG0Nl8+XNV3t42FWGLUR/6aHvua/TE1bn+uNT7MjF63
oVnuGfKTvhLe4g1vMMZNwQBHwg2GCGqim2dkkqAbN6OKP+GJ6/Qo2eThbHMrSdIL
SzxQuSny0wegNH/y+uKiEfcqIe58zkxMwZqSFaHnQB0x4CX941n5wItQLrrQQM1X
HV/tbRa7bFixCQzJVII+adBjULpqw/KbF21GpoBbzaSD1+2gaaZUkJQDAFmzbrqV
hJ2CQjXmi2ccJ1RSvhqgRaDdjrQW7H51AeM/fs45xWWrrdfu7Pm2VJX057oSxFje
u6BOeg38EuJaZ0i1TOBLWpmbuHAsxPk87CZOjYcbh/V6T/TUCf6bXzE0cw3V47CG
j3fAGZO2/nzK3ZRdvG+FO3jbnuTS0YJdLqmq+Bw5+SD/WV+8Ai2ftJ8NvcV1YW8B
SuhQAeLyYOT19az1EIvAImdXxidZiiHZupmCSjxR2sgjnxmBre/oo8a9J6krjYaV
5085S45FweWePQsQmGs7mDvsLL3itbZgA0jQNUMh2hwpVf3yQHoFme7lb/GHNBdi
XpUzLcr/O+meIpUP/tvDcccpkGQasMmOru/5CCTEHBHzKxftHAH/3fApag4F4EPm
DbUyr5Q4T2ZLDCE5akSFRMNjpK4ep4xsnik6mjE2R6RZSOUJo+4FYSVOdtIFWzgz
+DdSQRAFe8aag4yrJAaa+FMIkrO+6wIZvJEF7JZKBgLHhV0UqQxwy1LGK7IWpjLX
6yXfNdyTPJeBbvGbPBARZs2n/C5cnye2Tvrs3SUn7wjDstO48agjVad/wL5VQ5bn
A0yc3a49d7UwOId0zSVA5luXMpZkuRFsYYzHLdDrTjNd3NLM1Vt7UhAq6m2JPljM
iqeeeLfgSrIGgzHYYcafdo3UEPmBN1Z2tLU4dUvLWlcqQbpkYkh0xxN7Dc8TtQ1p
30pr+DMHbUknnjcWenQW4m+f5lHFtg2OODB3DiyNA9fQDYgjuUvsOyB3Z2e7134T
Htz3cPMiuj2JUT8B3ZgsMvK4jOsjZAhTDP8arpSUgO7jc7j74XaCfQ2tn47ylbtR
yo2gzqabLqGzWkpa3hETx1E4fE9dr2zWCl2aOG6VDVyIkA4pJSnDc38NTjqdz1OV
YAkv/wqTjr3xDx1v4aR8dNWdogvjXLXopiCbf3rlxTWd7LkPsOpzlfPKLoCYWxDa
YLxyGOMl8jbSJ0Oh7r/XKKMDA1SLggAY10VM6eFWpG0YbJBIWXRxonPVKKDFlsYx
I67+6pFSkEZFoDAKDNKA66ov6DfIlsgAMdw+dQLBt1RQsbxkzsyEkwJjiE5n9UNl
9KxirN5/NoGdltobHajIJZvFiGfKzBTiX2CpPOJJDz67ixapWA8tc67sd9KzB/yQ
PMOT6GLQK3G5UY1VGYZ/X6eOSFGPx9jKnGvZoaQ4jb/xsl90EhvqPCg5kTF3asGV
eunS1h3RCzAg5sSqUM3Qf1EDricP8vtmS+UUK/sJ25babyuKeWWWwbUv45diQT3z
NHFMuGXghqibvuXkuyKR+8eLs4Gg7nhOUCkws5oOWlUTo17wAl64opuKoBh05HbJ
uIXL0SCsvRHMexhdP4ghpmBa7e9BfxEUP6g33yS/glrJa47iFhKV0qftB9XCc8LR
dhZpfITKmvshbUlglgYNvAyrFWSOgv/m/+LOmA/cowlvOsdedVygOCdw4j6Fbio0
0SKs+EtXkST45yKPSg6sbplMHaoWZC8c+dQ8wFDirRwWnUN5huwDaQFQ5H8FopXY
t1IqIa4naDobsUFulBbERNcj47MXaS0JQ09Gqthk35gRbm+7JmWMsvuj3qhFeDLt
8gtpAuGuEcm3//45BuuNoQmsayRlXxTJb3vkc7xcuJENuJcH6JJTKLEFFkEyYAB4
I3TexpWIs6Lvd3CEgSh9KXYeRwEEiemeRCRUHWQJp3rpjNdiB9OLfGpX1ny/m1fU
a3Lf53h5zproH1y8m+V5+PIoYZIIz4X7kVWBgWbOm7NpHcw7Hs+5T/2eWRTAWt9i
0DYBHvBtID6NdUY1g0avMBVkTXdZPnxOnNlhBlDbY7CnhQKjSEUKoyEme8RtayyS
k7xJMNzKUSlEY8fQ+jT/tserb9IBlCMi1FQlg5N8j5jfTH7WIiVf9fYHSy1vvMMF
CuG/Gh5TvWAL8+iPLHr7WctvhDHP/3PD3BNfM2c/ygGdbbsZ8x09cse4S7WaOStD
cgJoivUTSstQNrxtuv7JrgR2iXNoS5mmqL6cW1h8H1/jAlnQ2ptH9E1YRPD15PRf
Wt1E6Pv3FlPNWkP7t4HZZWBWd5adMoXO0/ULzfRx7lc1cyhxFG1O4/+oETNMzX/4
dA6dNLVZRYw+J7+6Fj3rFib0yMGvDKl2j2BX2W9NPQWSoKU2S/pHkrvWnp53pngt
HyAhKeqzvvzHAY7PNXBe/gABL4IRpmacTtzExMjN5EFjfVwGYetjBjecoP1nraEQ
+PA2gweC9Ly+TkM+iMSridHqkdvaC6GZ/7+mb10M8ldQ5xVa6Y5yyVPZ6qsHC9aN
4x7Vg7Y1kKEnp6J2aop4QBDJ9Rd+qBfFKAHfVmwRLe7daxInMNNve7D/zdG813e0
J1udAbhm/NiBlko4EJxyuJ57gjcqTnHtSZRS15ggEqpSo7lxAApLoQsU6KVImQ+6
/dpiHbtknNyw92z9PHYxDke9D66b0NLE+ptBJ8kO2qzKqFrnxmfSkSu2zUYYrMlq
aCSRu3fhfndnm7Zj0mDWrtuqEEV9obykRMk1tv4g9OMmkh30LlTqygPno28QFmEr
fNkWARM+FAr2BobujdxJUA/EA7oHHBjvnP/Fs9rCxIlnR+obzCEs4k7ZfmJ+OaEl
h3+8CYS5LgIiQTmTSVHr/jQTJyPvLMkcJGrgkUGk69EkcKGJsday/5QKUqD5Mgfg
7YpxdlcbnX/jwJ3TxJcZa0V3VfiG1Gc953EBa2egVZGN556Ot8lJ1vQNNFFCC1s+
pRZkSAvCOcpGNbLqa/DOcUaFoJVJD052yN1vPAsoyHy8fy4y5/Jt9/AFyO5gkVy7
bn0SZL2PErfnyz77r93DbueQRW8Von3Cm3a0M6B/AuG+p+mUyPraMfmpSXEitLOs
fEhk9nQqDLpotCBhmtKPhsJHc3Rp5O4QltKh/U7R7QFn6qUmyXX1xyiKpqeH2dmr
GqEKJUomozeT2eEsWqYnHF8TPZcYBJLaeoxb5tXgfVRS/oml4sAzzBPScTAEGfwP
TM1/bkLsYzlsKueqgH1qhzxxHf3EYffEDPrxBDfTC5hzMCqL4M66udi6cgYI/6SK
TQlrxUhEKBA/zwNRurQDjUMmVMbTFDhlGgW04kymY5G6Dh66D31ay/LHEm/oJZO2
m39JCJ708IDbrKgjIBfoTTNubYOSs4cnhZ7CdAlFXq/zFDN2NKcUqpVmMlo3buNL
gxQRdIP+KirE3z18CMtRNyBUV9czcYH2feBfW8wtXXd7Z3Vz6+qj99a0d913V7F4
zOLZ4DwIiGVO5I3+eKYtMgqg1nmOSR1PF3SlGvAUNPJ2T9/s5DlGXeiIUMMLz2LB
nZ0Ai607rvX2aynHqFhCjx8ide5gyR0lwsV9kX5+aexmk9je7FEJ/yJImZmGpsT0
krePuYQKIa1Zuk6LFny0ACQ/5mQPsCxL4O6Ais57VfZdV2TMJYYgHbKuA9TLQTHq
le9SrZMZjzivYWG1WKofLmhn/okTkMb45Xh+BEs1ARJL0537z69glX+ihwfTKctI
PYqGdzesm2ieozMB0Vb+8Hor4ne0JuNXyGaBt770b9Y09Atdp8Cio6iZLLLIbKCg
Er+KWIx3QISW66q8BpV5mfL6xSawFiy16h67chPJAvcVK8UJJCySz+aR4eDCyQru
TXM3QBmYQik4ucNSuzN1im9oinOS/ncBcHRyP3W7HUu8VztyU3hLdq2zIuXTgMhg
2N9MEuQOK7XDlFj12aXHkEKl19XyPJYez7MJsI/rEyEp+fbw01ruLSriy/ONWNCb
VTdlqRRVo9XYpV9s5f0Yb8rG+HWGSSmFnHl2PeQlDcw5BpU0u82aHLz/Z66T8z2l
eR4gv9MMRGeIpBh4SBCLKSzE3TYrDzy4mwBwk9KfHeXgMoZWY0a0JDkv24/a717p
RIIHzWCDIctuWZ2ZmRH/VSX9HD+Qwt1x3WHaLhUeG9AIe3VPbPHsiYC97UulrZbc
9INfhgkvK0NRHDnZnqSYlX1RTdxrxOPuKrX9Z6G4dttaFO9Hj7GxmJPHhqFMOYbI
GoeDiqZr6ICmoryyOMZAJMWh7lsofubT0f3sPKrY0gJ4c1yFN+TmEhaTi52npkBM
culYd7zlzRVRx9xsA90Su5USu7uW7Xljzr5RNLEaXuqeRfOEXgpE5FI1fIMaE7JW
T4TcfA08sjgZ7h9EosLjvynzCPtvC0D3P2GvMx+LI6cj7t7WuPKIdS/MiOMMEY5N
j/9bThtC1tWfAAlCKE73aCyxQUZzHPpLiaAK6Qa1aOG1SHyKdPUiYrxQqBXqaL65
DuGQIpY3vtbLnjVxui0/jygmGUOXyb7kXKnjLYeQM8rg54Jm2FAwzMVj8N7iIlL/
iDIRmUQFzB4jsaAuiXEpfyC4lIHpAjM9v1oYGFnl6tDABYKzSAXqY2w5JIF+lL7X
dygHLqfGiQ4dgRbXzuaNfIaeIFEQGyBhgL53O4D6lvU88GuKokEvlKGUmmXY+X6U
Rf6oG+coJ029rJnurtZ7kzt65JrTqQpr0u7MoW8doyvso6b4YSiGc7j2ib4j6rDZ
+KIxkGlFKGMOLUn7fbJm8GPuIIKOL6QDNrqj4HU3Hkje46PRVIz2wQv/FJuPUq1v
uhRimNc/xaS94Xtm7vExO4hyiXwNQ5P5CQaImIzYhw9GnzuEBm6/z1qHSTHqDW6d
4ikvOuifrgy7h53L5emzeCmtVhhNChBEMZ3O7qTAFmApimKdZRxEx2apFC/wPtqd
gV2aYtR9D8pU83j2Q5xS71VTN7f7cEvkYzcF6aBimV9GZRwuBM7s0+LtNYB12W7D
E55M1FQYfFNabeqJ3uq0rPUlm3ebfkIZV9LBiKXyFLTV8LArS82SwumHO+Sh+sqR
FlOCYsaWmUK4AZYEfsiIA9GfY6jtGqaSl/DAZsfoI+SjgdgY5iTwEe31ZIO4JX5z
Ku3eQADAfvhRA0BmZdVGdfC6sTNyTVz7JyaYjiYk7VnNWN0sgIVnBXExBHxXUmd2
vlt73yKZT88n2O0WVQGWQ1pGPv+yelYm1RUQA+9hgyQMZhB3HHQpELjIrj8iT/VW
4EHjVbp4clyQbQqAu0VbKyRBG2V+HL71Yb3D/zi8pC4gufIFjcVq4jtwska7eGzs
eOq1eCyEWGAr8+EtEHWc96ZUVY/i3OGLP6hTr1n1RQAchqxyEr++IpV4v3De8h7+
GNqjoKfMfw7YvGO4jKmks4BRh1XYY6braEWQGnSDauyftmGDLA2NgzTroGH4GMeo
i01+v3eCUqlF2J2VoBzP/rjni1XtBWIXOqv+Qh4MjsgDGGV0OUekO/zx1VQRl6sY
AkvAFv7o+7i3FLhyEdPH05gW0AYMjPfixDntOmPCi8+JxOoQpQR1jFhzP/VPHeqA
dFQ69Cj+p8KRlOLz/5nsyuEEiV+KaoXhk4uo/h8Lwm4TDNYZ1njkK1hKEP+crB+A
MUOy/bXbPSd2OXbQeeZiOg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lcnE6JJxLWj5uaeF4hKs+U7cASX7WZbA4jP56LHzVkC6DkHvJbhlE056rf/C2atu
jPqdriP7h+xPSR+z9IH6/wVeO0/KGCuUuXL4hIWOY/frHhlqbTGloEfm8c/vTyxz
PiWF4yxquNdnglFA0c8mzbk/q3f9olgw24ULhYOu84v/HRe0lxsM14nSluRO9TVk
Ml8FSdqTu+Lmt2wtDbq4XqJpPwF2DmJLeUxifIC1AYc7KGKNaKe/BZ2gSt/HafQ9
71qGr3E+tZ5Nf5thzJdcyfHwjoNE98ADB7IpX3cnxnLUFkVlXMRZmM/gpHpfHOXL
I3w9IxOufhTb1nV9Y0kUgg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
Eaf6fcOjrwaqHFaKwbyrcZ9yyg9fBWWFhu6I4bDhBZV7sMBs8gn5B0/BbrLkHD8h
Aj/djJPfThe61oGS3mNUr7cHf6avPpr/L9iiTXqoSYbUlzTTW6eJGubOTuH8a46z
fEMlC7LbBVcz98bs6CBqENn87zrxn9ai14+f1afpCx/9O6kXXNdAy9B3k5BiAHXp
ko0fwxh40tvP87OOi9kbOsCnUKHF6PGIQKjbflgQi2Cn3lqPhmXiWtFr/G3Dq2Gq
noykGm1lkVt+woPlzTK8VLvAD8oeJ3lGDmqEndtyMIiDZqsUtZv7FS2bLaQATjRV
ywiv90DoYyWUyEr9QuYeCDq/X0lfJ6ZWZHurBPofhK5te8vVKyNqX5x/he5keuRK
wL6pzUEzd7Z9IOwCMEAgqXAvQ+c01Bftl1F4gc1+Gd0atBcecU2Zu2p/YtJ4iKBX
aa1/XkAF9awxagi02rsFb3CenX5ydm9+IYtDoR0gL4CNIIdjQZmzarFs3yOK+E40
Kyw4MuhzMX5OpoTcjm+Fy5aiRtmOlagquTJa5/eNXtQ3VFKnmXq1HIzGarc0QraF
OmzJNl84E310afsOR85hRNRUDRrhcSpffIoj4vGp3ZWr9y9SN9XeTuw++aNAiZ5F
eR3KxOR42m8bksk5kdTWZ/gxOrpr2ZIugcHAjkv5ALS1I7yqiTjgMxhlcj7rJlJu
QSm6BlKR4GCzXD1+NBji9uv5gnbRIMf2lpO4IXvKTXkBywo6YZKxS/yy7jL7BypH
2BZeUHCe/beJHFYbHM5qzAWSfOTxfLjF+d0l0cgqRIS8k00lQ3Y3s1UFcRwHbaqa
Gwe7Gyd0NJB7nn4pcyEhd4Gb1lNNpeEliXocqnBwvoAXXV+Dokw1vERRd6XmS1fx
cd1M3mDDpyv2v6Ep8HVbq4FZTdhE7qELMNXyRXLHdDa5xknvRMNViuxhlVucVzzv
qUcl+ak3i1CWssgbGpdxFTuy+BZTBGPE3jqmD5TSlujARPUuMmUlBnRKQFcIxmgF
za/31YMKeOLP1A2IOH5Gc822nONqQniggz5cYAsuGiAFqzmXPZIWbeO+j11ZIEbY
pNt8cYNyPGHOfC7OBQ4dAlSesOMGf7XORSmTV6xWnxiyc5/t/uDgg4kuwVQ5WsuU
ViQ8jOzCYk4xjfqziH6aXr8bXbAq4QT/aa8IBgs4YF1av4g31PNL2qOOiQ9Y6Uz2
hiCrhQkRB4BcjQHnFKWjcsUET1RToBF/DvNSsxZJtI8oFzKZRIOsFs4eIQVge3O+
o+QScRY67n40eBufSRbOpLW/eTHQp+MNnCormB+ygoIwh98gUKfkHhvxS7qVlGh0
UdAZ3fK0HwP4Xbj8z8t5iajhOtzkBS8CV4YQ0jNOFu8e/PIV2OaAt8pTaZaMIUen
/9NoICMTHzTCbIWsxGlNWfU9abN9Mtv3IUwdj1anEobjZsne9qw6NBXdG7vO0fxx
VbzAG1aDKW8J+CU/V75TtptAGE/Bhsgx840rSD8F0J9QMxBl8T9TYc7fM2IWD9CP
6FNiNqRmd1O48p5NI6cXU+6SZd8/b22257tC1lDlnbtsXpFEj5gu/Cux76FrDnax
yUI7M8Zn86iMSptko9ypM4dDUAkNUJpc3hEM7DbQS7SbXCvaXj7JtpXxUWVtca54
76aebPPqwUw8n3Sa+EncZNAQYHKMa/FHRoqcKxfQqIIZNClJ5WZ+M/dRL0wGB7SL
kTwNkd27OhUI5uIXF13uVB5Boz4458y0yTA056VArEl6/GU5ZmI0P0H12iDFBRYV
9mlzVT5j6m/4Pi9K/J7GjJo0DR76ADgRftbpO3hFJoJNkC6+nYDvnudeUMfKZ2uV
Vv4mlwd8hkdO4OCc3r3lg8tcquuMm/2IULuEpNNgzke2irYQLpVqZ1jL9ls7Dtu1
ZODalV0sOLFh7ODeKReQBj7SA+Z5MyRsr6TNieooVYzgaX6Jl5OqKk8hz4c4/inv
dDU8FuGIlRHfgLqFlYxJOXZx0xP51NP+0uzlTISuHydv762X39WSZZOQBWmZ6gFq
9JK6HehA9rijhLNarM9I0c+ycLJrjzEY0cbmI8RpWzbBL0Ri6dqGSAn3dNYWlvNC
N1j0RscQWGhTXnfh3PGf60EOThgd0h2qjkyld+JVk6Dt1ciz4Ytafstk5NxoXC/B
8Q74KjQ7x4v3hJlobUhm52hqDwSxTjYfnqMoY2yDWuy0krGCdQSbEFbvI8EIqdXQ
Wpmch13/shdt2sTkav+nd24lgmWvviAy3FxUdN7HUWb+8We6fTtRpuSquxNM4Vo0
duNFv2kBu6322rspN9Dsuvunn+3zEjSVy2pgyBn1VDPticljJyXOqYyPgXT95BwZ
xcDqfdZZ27Q+zAiXXpj0G6N3uxiMSjsDwO7G28Tufb7gTbwFoljPyVzelvD1JRx/
6gs1Wsb+Oz+m+72de2kRxuCOOlcm+MKy7NL5BeBgespN8Wd3TmdE4g/qFWSI/aYx
Kn7EUbeu5A2gk54Vkw0KZVYXCtqM7co/WJV89cyEqrXrMAr3bxM5Uw51h4dPhpr2
YCrJnl0STLTqAL0ex+8rjqQTvOdzcsKGhWtPS+7++mgYDmc4JEBdVXartemYsbk8
kymvfdr4vUfBDxmmRxE86ATqAZ+nqySfGwi1cBuw16Ggvh/tJO4E9zLka8/E9qX8
akAgZ3kgmT1icUmClomWuJDN+Uui/FmNjQisFVQg5FVxMs1LNqLtMNKduUrIGhek
htNReM5PkqJzDAQF9ij2Muz51y82lVg3+q7f+0t681me17GKvZaP6KvqLoP527G7
5ZbgBRpYeZFmsFmHfz5REch7qGf+Tyk3HjIqUAWbW+KXiisex/gR1CzP7DjgLUUe
/2cNRVO9tqYX+Age+lVIpzAqsrXHHixupaN+jGFngB6F+LL6swLjv8XMgT/9XRua
WuByyWqoOg45vixnIKAPTzTOi9ma6e735goSL/2XEss6noy75MjlChgxbIUPIvhK
k5+oq0UWBDIpQo2Z5NG00H4NdSBWeuDkqwD1TDWgg0HiQPjRyZOCTQHHBX9B0RnA
P7z7nsVwKkbQmKtFMoLAafEbFrDHkG1JNvxetJy3wPAeBecyyGvxXjtuisqVfKsw
zQxVnHxW9CalN22eoatkNzEDcI9kOQ03GSUHjjsUhMLfMDw0wNjW3yqF2qGpfzQz
Dz2k+vkaRO3n5WAvbBHl/3tZb0rWJVh5ZS/b8xJhn2cv1wLwlpMOx3X2Qi1vLpzT
AGJHnvLBI7VzwXwtgbWiblBspqaQtH3OrXRRjYASCzETyPf/sVmKFV5Saq1RWXyC
PNuLW78ZFPTGOw61w0QpkQPylmGfJ/xH72aPY3m10G5vJFUmxJr1UJAOY4c0luG5
3tE3sG3Skr2I+Eg2ORtT8S3ca0o/oBXyrKkf3ZpldR0qli3g3rkbudVZ6AtPggH/
VDHP0jsg+WSepPLq8UcXFo+Ig4buQu06uziSGSMPpOslk2GIviHZ8t8VgYrrwauS
l+LL++F/OpTwkalNyNxsZHdKGzRxTZEAkRHZm4HBmw24mICcrT5YBlmGHBSQETRU
32TWU0VXWLGQyH2uU8TiebrZ7Oc/sSsp2O9iW3XzVsr7u6kEF6EKtDGy0R/YsXgL
nZLm4eLNZNxKR4hDYiakEowIZTVY7MVfQV5hvmbImWan07af0xK2bmx/x7UWARfi
AemGhh9AIe6EsmJUhhudTpIVheC6mY9N7rxN6HYwKrGamjeJzS3Rz5pfZTQfk85z
Wzid27dj6qZaOIFU9zEfU5xExhHr1YBArpsjQkEeGbyPuiJ3gYaCkP+XK4wfm4sK
Vqs4daaj7pk+ffNrGXRWAdBKe+uzbNccCaUYpa0vu5dZqdkBr93NPTgfGIVPw2SN
lQ1XB4ZK7e62uHmJOwV3YmsFtm8DcKqDmt2UcSOxSc2AMutQ3zcGDDK1EJ7sijfc
Jv7IkV6KTXl20QM+gj76db1xfoYG3II0eBw6OCOGhhnXfdGih32uZdNdRrTuy1Dj
JtR3prpSKqsr5xszfSSqMZ1JF+Zh/DYq4wGswDfqHchMZQGQsg/32udiBP6kDsw/
kbCfnthPf6o0stNF6+QJjTzEDijo5VIPAziNbR0xOvCFxWG/EX6qBoPD17S9nvCf
X1xrR95rqcmvXGYfeBwR+RPpy19xhS3YHd0sd/5hKW45Jf29wviJ4ZriUxagOhd9
iN9EHU77iaP4YOVkZeoifL/7KXfrVzjg6V6G4tgZcYROlnoVWoYcb9AEinessza+
OoOTM6fYz8rvk9sH/kKufgq5Dqbmefn1mLFVxHaIAnDcOKlck3UwtjTsZy7k+vx4
dj9POqTcWOg10KKME+HvTO0qgx+obL1aTcMYtBE7Oth6PgQ2ZJYxDt0jmKXYjdfO
5uCs03tyg4y3cpju6Ml/13Gs/+PiHNrOWjGdmlGykTV4UkHjoriXCVry/7v+xYx8
+Gm1MsewXSJyzEPlwLcykwWvVXOIL5u5Xnfkm53LjgFxjateGLrFnAz/R5+BWz/X
sxAY4qn5diMNhziBksXrjRISZ1b1coWEj8V0JDEnnmRYGGqxyFnfhe/2v+27cDFN
x5H8QRop1tqgDI8e8kLxa44mIHykyyg9XBzDx+qTyWJjNjkEWt6ZD2VLHZFeNc2j
mIVAMH82waw+HBGU4+6aZ0XSC1k6oPjClhLtkzl1UNsICZS12hcOW4xtz0lP3Asg
Sj0RG3CVGyQ/iK3YSzczOVX+0x3pEDsX9ghrkaB2WWNSBQ2kKJuaDm3zkjxiGRiK
hxsCfCi3aUKQAfoy6XKbjy4HPcKaADCgnpVhYYgF0y66aSoMGLgvgSwGwAg1sDU+
jVw0Vn18aOpT0v5yqe65RS9cxZihPzqkVr4mCZHXCWRnn/kLEox/ue9QziTBr7dA
0lRSwNldI+diRNV+AnrI38VPleaCAyu5Ds8se3v+4UbTHdh0TJECCjeVlV7mQuuN
2o124U0h4sn6N7OgBgFcVWjFLzK6Ude7Rqzim4zXnmdnD64JEpgVyMFejg23BO/X
UNvSDwJrV683H+AkrREWPlpXFOlQFIWGhPTb5Qanl+afhh0BA5VSrlzkVtMMDy/e
9zhEv3ShfLxZSSQGiYucA/LFK68aFtmeqVu7rDOTzHQL5rFoW6IrRMi5OELDzyTe
J4mrKaOdQFgjCmTbDnlQfkwc5IRSy9xxOkYx3lzC1lhHt/wZoYuAJzvq4e4IVqeK
WIkWZ3D44uQT6RjbrONVYFp5p0uCX649Co2BvkOfsVAl9XfrKpC3PAZPxdtvlzUz
Yu+N/7715cHh/EfOcShpAtEpdYG5V1lrtLOlTHklLpB4r1GwRTdCO5DUniesLIw/
B4iEFWN8okSQHIv6ROeom0X567ZcJEKLOQ8jScVGbhkvfxacA3WO84g4swxe63gV
oIAI0oWVmKwf1sNBvyiBb9MxgUtSDVtF7RqmtRs4jySxEP+JSQE3UocuhqSo5n1A
UqASHJn/8dKCJrTXqslau53v0f5I+aPXfazNdvcDwje9k0YR+Ttc2jGiCnkoWbs/
dmeIldqA+muRpbQ26K50TnBoIF4AFXG8GXa5R4gK0ksQfzYiGM5EEDY0EbV422Y/
5htguW5dV65X+qhUm9Fy3MOtO3m4kfLKK4lKILfGQwNp5rsMtVnLxydg6YszsfTA
1NAnYxV8c2+lgHY7Z13FndOXEkc9FXAD0a1I4rwiroe84+aG0ltVCy60oiOqxO2P
BevtYcgJ0ECmWfSK9Dx8l6D/fSKY5T/wziY1sCpgvM3eZ9eS4laRJzBcPY9ICg5D
GTiKsE7USwF8Bx9OEscx5H+YdzMVSAIKAd7B9uTACTBe4KyzGmfiqzVhh5/qoyyj
XwzwKFo6kNawiSsWI2gUQdWF5x5V4XPzHZ8gEe5vz4/ysnXakdnOT8ZoCiDUVlsn
1huFhmmqAZazKOj6bBEsRYUL4P+JhkK60kqxVtIyXpjEzj81wMjqqF4F1fjuyHhA
D82QIkTK/x7kqjDXO3ikRdNgCUfpneiqXIc+vKEpRNwCjSZgAm4ML+wjLcMA0AbV
b3lsEwpa78H38ctsGA7eE9GCIY7cWyvlhmgeczzvSNnaW2BVn3TX70v6IJALVM0c
2RvIFn8D6/o5tgwHwfqfa1Azi5rSlr9qqnI/dQvL5y1m8VxhtEmmxm18X/icYTFJ
gxARVC1x1r3Rlc06O5RU8A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BWx0iCnMaaqEllq6KjbfeiaHuAESxgz+ua5qtX63SXjFSCMbocQEjPouOjnXnOs4
KF9Ibva6eOdkMVArD+NSjrvPtxSg/E/B8e9bn+eod+a2GpifcpazpqoRVVbg1soW
LCVGWD+Z0JKDd99cE+BX7GrjH7Lf77ce3so4fWYNvKoL/IfkuHUf5BpW+vUckJrr
A6xoYghukp4s7MWQs24BIS1Bgn0/+tjjbvATBdOlWqqoIV49SSGy7oRpsJRAKXX6
DsDCB1qGYSZ2WcCmeU8CW6CQU/Iqrh8P1TXfbbUCL9Fp0ZHwTgnl2SRsu7Oi1DUv
iYjtMNW5I8J3nOEgycQN/w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11552 )
`pragma protect data_block
VTXcqjDX1KTzVFrSGGBlCRKnrNGRkDBJrOSZU9pC0csfiW+ssdnAPUQ/TTnno1V3
2aCvewFk6QXhtKEt/iTQ1+4oUTnEaPiALJnkIUB4vsUAVEuyp7r0uwUP8ImmdFU9
Wj0PKwn0zt4724pBFsfrgbF/S0QUdKpBfrhYBSCE15MT2zK1erB/o7ZKCozlwQEu
jrKUPkErYiL4OiAht0ZTwnU7tPZxnapSlPmoEqDCPucAt3FkAdBNU1N09lW1THM8
uRenGdqiPKAmHeo9cmEyDXv45gr4BTpipBZE4gfZZ9nqfqz2f7O/UsOoOyf4Wilk
EqFP5cEG0BPogDUs89lBfZvqha/xutf9orkgWkY3d2hmH//pTQTEy5HWUWisua4s
1wueq2U9MD3SMj8QQlURvwMnlTgkVQkuOIDpVHm3eESgGYXCwuk5n1ruD2DMzcA5
sKsvjdJw0MtAn15o5TscykIiyJnYj15e1iedRquNHErUPUrE8ajiq0gC2VYr9hus
lZfVcEsyrdF1XSFqamZE1cslwiYor3cnSaYF92BbrHNVexEqPNTCtGZCTuf1INDn
w+XecHgD/4ZVdiPPjKBunnHIHpL9PnZQmHR23e7sWcq3blK68AQPswIIjn+rFRlo
gg+uVoMiIDSML0FpfEKBG2pHp5cBn+JdzE3yJqiiLvBakr0h/O1rBxrPhCrtLRW/
xRQFBVFCxmLjzw9mUUJpaHOja+KLToGXjBsY5RuDbmcEt5YBxpjoOYYlvqfnkE5B
AGZfBFfDsl16ana5kYcfX5u7CZZNqtMLs5BnTkbS4H1g0njrGgW5tMJrPUSt5I4y
WJcbtRFMGWy/RAqDVBQEQHJb+/N21wojgokBEUbDESBPEXfwzfxzdrAwLRQI+tzM
8w2tscOU5ud2jsOO+Uu6E5OMauAfooh33r5Mw0Cuc+dxSv3p58XjDVVZVbcjDb6X
fPvFE6FzDnfgHaIft9uOkPFcUbcaSpfaTybNKsuoqpQEoo5Xp4FAcH7tuyZN7kng
IfrxuqsnVS58SNV1YvFY6e/yx6hIEQ0adOv7Vd9JpClnHcl1a1kjZHznbMBEljrc
aFIgWikZBzz5A7eaJvxhvBoUoKtv6N5ARady0nlmday8dc2GRAStdOdkgvdaqk+7
lz7CJrJUBgbGNl0Safkxak3kS0sLSetRq7Mkd+EU/l28z1BPhBld7patv6MiRnSH
xaDaQSJdi5bNIK37VTn8h58fGY0s5IRUoR9JUSL0ptDz7zzUIES+DvA87v3bVDDG
azhrarakcDg4FsRvq453nVWz3F/8cvK2eOXU5oQ8wf/HboajZlr9u8mrscx1AEyw
EYa3glL6Dbr7xm98+shp35TtBAcQGcfsnsNs0zErY2R+W5ylQvDuSkRzjrzsAW1d
UHzjlJ/lO1O+yCcUnv1EdLhjx83e0+5nD9YuP9u2oBFUJqOezNaqV4uXgz0UFXIf
ePvUDYWw+kuY83pLdeFBOLzHzetuAWIi4d93ZkGg/2w/5e9Ok0nCE8gc/gbfvH3z
1uEMKRdHuII4aLv5v/JRj48zzhrm6s+Ae++gGCiOAI/nP5BT29p3ooYDpXU+D8rv
Iwn33UKcaq4LZQrmMBA7bK81EUwfgrVdEzPdGqdkICTlifC8AZxhrxuDGgzBxP4U
Id4Hd4hai4JAgkVt92DCa2GPPYUNQBXyVhkB5Usb7oUGETg9RiRTHkoT06QCIBt1
2Rc12ZGmVmWSC8bVEIdLQAgJBWC0huyk3icJ2qSpnbbkfisbXuEtLrVrmkKMxit9
NZbY3z5AX93gzNkCL4QRh2WaMGnhvbWhtBLGlxPaBF8f8N7jsvOnxV2x3KjOKcCg
ValzlK2/m8Js/ftpPl4XAcVzAcew0tjONsSbup1KC+8Wg/JdjFjf7NFEtMwpuX0u
PV+2qNWxp5mndKAhpvACVwbpiOezsRKEJo3q6DPpHvGSENpLokzSiIIq6PBNdd8G
S0CH7UknRRfC8By8YsrO90PgvGVHjAuq3lxVTHJJjW5NV7+mIlI7v5R2jEcK07cC
4OEq1JPAVrnQwgc12xYXQAM0jeYrR8iqIj11TNJD1tiki0lCAtFxKDublFh/YmEY
EGu8dRWT7e4xMHzrzzm13fk0oyOQPNvg2QgV5M1PF1DqrUAvaODGaZFBsnmKojhb
hsjfvdz6CUOoauky5ZvkxosrsHANE329JIZo7YE71C6DIUGigFQcB2DHvWVZRpx4
GDsbZbRsJxPmVlNoSobZ+0TqSp+Oe3foNAVgeJ5SlvhEvJR9qvU6817PHzK/C4QW
UheAFhPhQxncP8fGXJ4le5D60Vl0VzIRQW2Cf5k3CuXkGHqqz+iJFiwNUJOJMaRk
m+MhIZzCrr2/4T+hAxpL5ZcX3Bu9tuVnxns4OMABt2Ov+tle3K1ItNf6X82er+sk
NrkCWhFUZ5211JYQiLeskIbCSjQ5gShdhqtAyjQiv+wYFi7TukyTQZ9exsRssIkA
cObEX3WGKOpac4xp09Ogtk5GXN52Ctxpaj5Iy76XQIcEsPLE7nonMXxTMiRisnkz
giSYVrCK/9VpsWsZaiPmXyIGtjAQ7TMtcBanXMaoeGtDIpaFEFY/mt5Hmm2RuGuZ
2+9YE94h4kYXQ/bjgw4oTbyCXJ606qoT8Fq49s2Nyr1BpYyGrePc/m1B8XeH4H8u
shgIE3rW7vWRMGZbzfsdtMDX/Y2UjxdqTwZo3LeAfeeyorRptJhAbSyN1l98rbfm
63Qug+0fMwJ7fysCd9cHVKDx72qWy0V0qM9ocWim+qBfXWl+Y4BpvrIjgXoBJ5wh
SyjyZhcuiBb3XlSls3+2nJyqLkXdCAA1cWnNlpDND4JH3JN2WgF5yGzqDU18Z6+g
yys5hAgjQKD4u0SQxMz8qg5tz25d1Z7rb6lEXqFI39WZhSf0q8ykJXBBsAmyBBgx
m2HKPbgZLFzkm2ouI4R/1lR+tk9vDcP1xDw+ynvcx2FlpWeJLBVvQWScr+Ud5RW7
lKmWzV2HisGnYBQRLRPowS2Ad6N46JRTgPcLVrDwycuFN/FJKgrU9sscZSOTN9bW
VHIboJpxCQRMnu3BaANeZNwY8OL8mbn2PYkiSsxdi4gNX4YzB7Sem4SoKmYXpygU
+TMXH9FiKGXgCU63qGoAzwMlnOR7W+Vr4LIjF61N77zSyJTuMxl2ZS6MkOv5xszr
6a9MPhXXFuv3i2byayC989aVQ2a7rMykA4JHlof2NPoobP5XUOLCWQQEKWMiUuBd
UMBdv3Gjj6ibP0gfMFYNHNWXAMUEcr8N04RrTY05NcfT8uF2LMs93cozxKiXnXhc
AdYkpvIE97XDUvg2evSYMykc9LDaHokLBadmqUno7Y3GaB7hsxAO3237gP+bUEnl
ZUcAhJGQYLHsBEkpYfU/hVFQjBN97ZGUXKpDHSw2OSN9d78CkEue7KZ46FNR8c/P
AQQlHTC7S7W0+d6oRFPQ6mtVifx7Bl4Flbdt56o+JdPqSfdtwInSCJzsZ6QhB7iI
hpkfSVKAKEGVKZju2DmiglIw3Tsi8UbFgFYR2x3Ov2Xv5RXI7loadOjBb7W6Gwle
lOvj1eVD8xIY2pzNSOUBeZj9/i5VQy9Hc3j0O+2JnxSheB6KfUV3SVvfH/XeK7P7
0uRQe04Bew2IyraAcSuHCRMj4IhsY1D+5ANOOplDWUXW8Jhi/Dr3Kmq9i4G9SW/N
r4XREXKbtSVkwFsN4dOdxi3QOEZl7HcC5THLEU8wwZwXsKbA44ea3DaLTiL7YTin
vTBp6wSEt2tHn5RuxukzlutA377tYfpthEXYZ4WPzdXIROF5spQxh22xzS6v9pfQ
zVpjk7t5vD9bGKvplBrE+Zr4mq+XXjyazm8e997KRAPlE/Te/xj2Dgp/ff7vbuzb
jNfCm7Mn+xw/MCDktm+XN16LI8Uq8BER4hwFU/fvJqtHs5akUxayCMLHveZDVeTV
h3fIOZ1pi293LwzL9WA/bTFqPwZA5ALeYfeN3hJads4xxD2QLWLtkNsxS28yFfUH
UuLpX0xTpb5q9a6wRCHbzVbrJ4wvH6ejy0HYBYWRh/FbVgrLnPbsO2kGNjOdpi0s
cXFgUYu+P+/l5zkR+8Sr1Qwbvp6dkTDi9L+rbNRiRvpCItpZfMLVFuUhZ/K9Jdk0
lDoa0srwGfhyObhlhiXEnVCHrecq2osOS6GqzqnbMHsc+sDw6T+2z6CxKLSIYZFX
LocOHCSdsus5Wh+fq1pTAwVwkhtHluqkE+ZAQY5XBPPpB9+CpCIAGo2GemeLm1Rw
OTOiz9suJ6c4nII7z+zSY6FOA90NDCX749QMUr6wcrniWj2C2B2zaTLM0EWdZfV8
PXqxT9uTh/3dtCS1Ejm1z4sWShpv2rnJe3C4/PNsezJQpn4C5xMNhrNBz5SsXkEs
kgOM0QVLTpxAQHpVu8c8CUwb5BEu332/aU3kMx+wl/OXew2N8X+tzqXNQSsIfJlH
c33ZA/u3/Y+9+8FCvxf5BAkGc+VpOVFtguDUxne0mfjDlgIOrzMo8d9ckxtLQ5P/
NS0PZ/yfIElY6792U+T/kHnotY+WvhN7/38wGvjDXR3I3zLJ3x5vgSgYLP8Ng1S2
9k9Z0QZcS0B0lAzUgwVR7BlhmTClplfzNOSw7Fr9hOj21tbZagVerz3KWu6DD/4f
tu9hUyMAvQMbSSbA8YnT/5N4fvFoSPVOqzHNuKCvv5A/FhMeqOsOXNX0bukv6Oe/
veOSSPuLmeH/ygKe73yddELcapzzFMhCk35AkDtuuWRSaebDwyiH/OfSrqgy/pjA
DnlJl1Xx6xjbkuKhyk8M3HbBINURMcy1NtwXkQdgMF+XP9TiKB+mtIhVdmJoELut
PnDCanpqNl2+EUi+8xQ6bMh6J0St9oSagXl21I1Ttm66khef6nt2xjjHpNmsLP/w
o8J2a1Tj/CVZhqkj22L+ZeLInBTTiK93b4Mq09b0VLhOpMwmFspOcguGjNcdcxeD
ve7552snSjsBFNKVfUbbzmDyH+7j1kKgCSdkdGvxAjXqNJCOZThop4BTX07aXsKx
Gmce33q0eTF8CqA1FLuMbT+NFLBPvxpsKIjHXCEUybys6xxPDRPFL6yzCuP0zAZs
YYk78TmhsSFmdQSbXGpUkgKf7vcNSHt93TRhRd+1hgSs1aMh+y5dNy4nwUwO8sMF
ebEgvjVNO3IG0HP/5MeL5snD+q3+xPyxAXL+DKt3k/lqCxRhLhk1FkAHvDfE5qis
WZur578PccxZcp8hrEQFi2wsntUrR8MXMW6EAUrQly4XEcZyXF7D4vTzL1IMDg+k
nFPrVsl2nX+jgz4Rf7F3Cu80TaZYK1dZj+KtbKmh1ZJyPPiyIfZubDLBf4ir/c9V
pLNucQGTyWpJ5V8Zhrc55VPfKAy+tkcMo8pKEEDd88MgfavAIgl4Jn1h5BdSt+Vw
p64s0/4gPgAAnwGCN9jK9UZwywE/ZgEDCdv8h/dV1Zul5ey9UNKWwI7kaMa7jcBC
6rsxzezclM2tZm8D7nkefHQk1ou/JN5c+CyasYOTRxiIJlpCBuQxcNlunAbmOMlf
yRyqVo3e0P3duq6fMxC/g9qy7Ly8Ha+K4DT+Gg83791cm3blJKgkPrIcVODSuqf6
GYLCrRmv4WYIC/ch+QwVsCaRLSg3Wg15MeNtp3xMTMhYxnDsYdcnVwUac5X0UDum
e9bueiKti7814961lQ0mH8Js4r+l34d0wl5J2ymEc3wlnZM/QRe/KxzThK24cWK8
oE1p9zT3dMYYuD/Ry+iZ+SPC/S8jqrNL27gd4wSGFdZzed8wPOizPta/D9TL+4AU
xr+F80Z4sxAMAK47/1wrP9AxtxqRHJkATmRkDrB5d9BO3ZmCrwePvhbRFHEtQ/W+
Zbcfck+jBzdaqW974x6s6+ajDEW/gZjZiP1XAYsQ+pIPiUguo9I+j/iL2msv+HBe
VUpufsYGIF4G9gm0tW3TquiR1n/EI1woz5G/GhNj3ltk+cYo1DBvPwvUq+Y9pb0a
EiBTWrNfyQG9i5U4pQNaFCec6K+9wDe2QSQeHLmvk7WOtyidTyEgi1q29fX4NTH4
glNqnvS10bWe5dsBRHKr1+JhCAjFxc0eKuHN0VNLLaRZV+WPEvPS2OuwNSnFutWp
rl5fixLWNV9DC/EQna3Owojh6g5OXA03N52KJm5LqLQDmizCdCO4G0tQIeHMolJL
SHUUtX37b+BlnP/P2Tot/PDqdzcBcCKL5JxBhoifXTasXokdUZ5sS3EMOTjrKDoc
wCRdQhEAfUZ0jUiGDcCeJOtkgRhiuQunMPbOn24RMIqyamQgQqiTCnV+nNisHcfb
PuPoHgwcpPq/x7EYaLZwnddeOkRaAYeGbEXGCzUQ6siXLrp8oljqVcub4O9/OPch
fE3hXohW2zfrzoz3vBR6A/I3alxM0ocM524SVnJe6ilWEWhDSRim+YWYUUqWu1f6
N93zcDWyp8Roc4nEcX+sBwQBFQBpZ4KnghKTYp6nizc2mtdngPhzYAkjWT1TiKGa
SM+boLtQk3++fKyL1EU+GQVJLmMLnpqj/PfVe4NT6zhUqMsz7nk/eV0JIe7UUTuR
GM0z77I6OAo7LCPa6xhbAVSQSqahYk8binrBDB2TtCeOxSzwqmJTvcOWAVFu0xVC
XZuqLLPXd0bjXpwmjL/atL8awq5/P+N8SCEl1C+W+/OA794sNzahbwg4VKUi17ac
maxdHwC3fpEy80yIT4eiGIVHhPQfezXwxEowN981qOosmioeP5a3TSrSKlzBD9f2
/w1nQQ07fA0ZsysIlcBgVdwO6dA5gqn5lGjfer9rid4+g9i841Y8OK6ykCHLM8jh
+QsVmcVCTsp6r1Sb0HN3GzRHLD67RTwTCV7g6VJPwwAOwsdZ9oSVms5ypoKU0W3H
WwRg5DNCHy18VGz158BnBBW73zfj5twI/Ulj2KK3mFA5p1vWAd4pXLX3RCif0UWn
KGAkgfNL5njtklGy6kEL/0Qc5Oe00LbBwgUPyQOV4XqfJSTA0HnpRwfLrfNLhokx
3zs7kl3OIoxnqUssbSbRXFAv7MBH2aH1C7Ka/eZof74Jl4I/kr0/Q1YWBF1YgOeH
EhCB/5YwNykkGfrxy/5ZrswE65i99DUco69AHzrVFXOsw2l6Mqvkbs3bV3dbfr4b
SqHxjDb0g5UliGysrzyKL4UwUIw/I9CTxZIFo3v+IC5EUjYBxNr1cO8nAjIV2pkS
xoKl9HXoE44xf3KCqYhdpcxwiBLr98+c7h+LzS6ufQllR4RvOCPdSS9iSESVYV8k
lL29V9MVJJsBEyz2TE+VF6E6RM7ube2eAYn1pFvwMrQYdShII17Qn/aLPx6uyoUb
sBg+yY1y8KeO5nWLbJDRgEoPnJ2cL5kviWGyJ4YvlmT0whPiysGcGsMEjLonACSC
Rpxvcw7/q5KLEI5VYhz9z6D9D1zH6CFyI9X/A2FrbDgqvVwqgJZWi9Fk3zF1Ww0v
/MQdlszKSAlTTx80L/IHPcJCa67rtYpWdrjBCj6MQsocuckVdP4aHSF66C8R+uY9
/r/C5v6TdfMpRbOB7nX5CZDC95VqPTwvu1FuLiu1MyY1bbX6Z2+YoIxCkS4TQwpB
e0H6mHVyxF/lp5rAaKxZWmOaXSLMeuBPG272Tr9x8hZ/gKbom6AvkkSYjy50rHrq
cmnm+/dFCyI33qRiJolu7xql0d2SSDgSvQ1irxcKS49tSRWu16wQp28R4djaIOCA
JZYlFCtk9hYIxnglwUJ6PbxJfmbHf63L82SGytGWX9E+lA0rXJ3JQLj1Pahk86GO
RPwSwR52lrkD9Vs8CuVd8VG2+sBp04TpnSH1ZXAVLUrrF6Kt0EttHA+vGygo6FQH
Wr6BTL5t99KLK6IGxG0PrLyfz8Rf+6qkbXrsErcaurXy8y8SCCWtuSqgMgkWQ53S
TS2PgbP1vEfSl4sfHl2F54S2LgLeEAX38Rz/BkkXrDdekVcGdR57gb2RHYR5T+8b
FhuW8mvfbm9UIg713Knu/mUAPxidqYAHnhjFHa4Uj105FqbN9xOiFCZIATyIWOfB
/nSvFfXetYU6m46HtKYG5W65NNy/fqo/1+RAE4JJW0Tfi76eNbggBOymxxuFraaB
qJ74uQ0qFeSXrrMngvXz05g7yaGvv6AMmP3BX6XtFdvN/JWoGGhHQ397EtDJfuLE
meya9GZGpot/rTMRnq+ncVmOMV95d9uPXNTIXelDkPIIAXUcE3SzSH9cNJcnDw9x
LDKCv5mG2ukL+avVjLtv/1JQE7ElR1vbLNmkdb/zcqCmt/wLXQXiW081PI1hZ19k
SahVqRYRGR4sZt+oVKq+sprOyeLuEDWGVvd9DY95Va5PGa+zzNT9sF5R9Gv+uElM
a0LoCK01Ne7qYXJ+cUYtOoxMpbxfPwURCnxBsvBf/MLM1Z1o8v2Upplsy3qY1cBf
9XVzM1qq64gcMHMT16qSBIVrxKToEs8uBd87Bbhcf+Nz/bjM0BOUewqhq3qfTVaa
VavlFGRLHo0KoYmGUg+La0eCDIiUMByDOrQBMOm2A4QY8blkGRM5K2cHeVeyCJFD
oH4Mb8+65Eejxx0Ph4POiiOkTj8vp8mFRQ1JKNFtLH9oFfKXTA6es1MoMv23wLSv
h6JFQRYJjfl0yf835cVfoAKH1y3jxL7+s4fZo/c2qFjEr1Pr8vL2RSt7wly37yVd
DsUNa3sUf+RPfeOaZYZaIIufMfWb2LkvYSK42hDxgsg4rcToxBnPrrHBRWI60Uyt
Uy3Et1ja9DdQ8Ax7BjkQmelUITAGPFOopnFZEuCWYR3iQhqXK7P6k6Us3P7H9q5M
UDnLe114HNU8IOEqHdMabRSQozxZYxrj2PHycEICGPV/TOsP+LUrhTroZelv8DrJ
C/4JDutB1WEg7PEjUDizF4ENTWmWD+vXM0G5CKCzOoJHMDeWlkGzihSJmRqQ5TNz
OwgRnNc+ROYpz7pH6N86Ro5xJ9aeoBBf6wJHW9sut7/AHRKbz1VfIfBRzVtrSDyL
gQkwRxbh89d9/+7JYw2xmh0YGf2cs03w+RpDl/7Yk92J1IYRXt7US7LCtt6h7pmO
8eI7XOrFAA/bwsP8uzLrwl4EJmPJt0CRep8UnMAFCgDxIOEJTdwzNq4rwt558ge5
Bpo6f7Cjuodbglwhee9hNmv2RrQqdDaVF6hWk8rWcfWkiT1F6aUwYxkhplTIC46M
IQgBcmUoG4n4R9EaGiQxhsSNo/YbqKwdfGxqjZqes63pDxpyyCVbNW9Cl/bb6Op5
xVXNheqoEujlBj4ZzMbC42F5OCCET/quLBiYqds+Qiawqo7zl1Jjm0XJFmgR9/7m
KJOKFaX5v0ECPCgpNCwHHqPwLnFwIqtWkh7P4EoVKdEKHh/+QavcmjOp2uKTKwIq
xdBkz4kziAEyj7WFpNp+i71YUoF4NXibRvrduxQw5yuqXsffar5jEQHu48ngrGjC
XRPkAo5+hjeACIHC6UwzSxtpR65+/+MvbgjPjGy8UR+GG6Bj7vDpYIP3owhS0IXg
X23ka1uVqc4z35IJhtgwHJA0gKFVL3AmwhVpRH/cEncWMFJ26yUN730gz/4yWo5x
3OwStJSABk5Yn5OKP0MFnDjBKo7c9gmr7hrdGkxyy8HSB8vRimgIBBIPJ9gy/xVZ
Tl7BY4lxc69TCO1c33XEW1TKZG/9oppIHFQ8Xtl52jlZV/IKjGH4qvcMtPPRvpTw
iX6LMtHvwlJ1YRMAnSTyzYFTm5e3WNC3K1TcqaWPhAebC8yenIiDuVZNZz3YmZCw
wE7Ms01JPZEAcbbJPuikiyf6lX3eAPfaUjFSrPEi+0Kf7uVqZfuy56CnbZIsk+pn
Dd7bP6jK+RyRzBerz9oKIpirP9p/rdHE/9zrtRMDcSuY2Q0wA0pUH5dRdiJ3HHiY
3Umto/8VpyZV2exPTqI7WWzxPapZAgYFaURqTV1lhKFdnnrh3XUUxgzEuUq816KD
B6lhHe5iRt8eN5gpQbyJJ60oBaVH5BQn/OHllrtW4zacMtd2nP3dWI49GofFcwDY
lnlQaBLK56oXyR3qamITz/T13rVxBTXU55FFaEfCO3eUPanfNAiLonxyX+9+S2HF
GBuIx31yxM07pezO+tB+In/Tmuo15VAmqsF69ZEdfM2f12omhbKeXIVglR5cM1uu
oHNvHUXddsfJy6B3aSRSccLwExY7M3B9EXkCPuXuhPYr70i3mZLv3wPAZydymu0m
do2M7q/hTrNBjryqlzPo9W1HYJ2sfkdE+vkhrgqvxC+gvTOF37JPcIE4o5Wopvj6
5ISMX+Q5FHQaU9QDVN69p69PvTe7/LrpcEK/PMMJKdc79d+q3fxO0kZHF3a/0yQV
0keOC40EzSMxbmNRPirMlDam3PIDy2HbHZqTkMuBxZ2vGLIFQWjwUB5g/AIemf8T
/VDkJ3liPxdW/MAB3eC5vXJgrDTV8OpqIof3D5M2qIXAWVGwpP0vXmFDsdXTQPzw
TxDZoSksie6S5P5+raQpy4jqsSJziUYeD2ZGq1gSKVIUzAAGrke8pvfAu0nrDzzW
avFa1XfO+pNKnlqXwfoXGTaO7tSCjxeq3CJ4Bn1mL2cW0PaBP9Y++22UDYCU6Jvh
lY5qP+SVf/2n0vmazjAh9suzX36AmRyOWXBYSXA3sSf2RCKdi9vyOcz8nehbun1Q
pU5ubZ4KwKHrBN53VtGhJJKQwNLTl1iQ9DceIsyWyZl3jPxWwuE+Yp+BQE9JDzex
ui8XjlAn+QihDom+utos8Jo56wzO0jha8hBy+wMrUeDI7z3u/cgkqYDXigFSDJUk
vzBakfY9rWT1J6S4FmPLHSmt+2HxcrCOPF4s48WmXCexTabiv83sRu0VqQmirE2Q
vc4kqCP8lL6cCvkzWPbQO0mEZUDHtHqK2IlA04IoYNf6LbxyVUtOevnLuVgU/KQt
3PxXYqs+IHk73hliLUQpwDrxJ29ICviV/rvDS+8soXOZAuIKylkELAspzqBs3c35
fB2s9TMsAqNawNmdzj5a/IMMBlvMl/oBwgjzphPT8rZ2RtbaKmcqgIg2zNU/0sGM
YAxIpmH30yq4SxpMjFLogFYSIHElMqo4W9yqnbXUKUbSt0ddk3o0IBJLTZe2tVo8
n0RH40INYHSbm1lRSWVIB+aUQAmUtWbQ0/cPoCLFqSiPVd789UQjC7g0reu0HPVG
5cE6+i2fz8+Ph4DYgqu7zaDnZdXFnsZlQyHDLwTnUodsUWFrQ7lpz7t1+NKoKzZb
7XcKCStcziTMQEK1TmoN6amhwIW3eNMm1r5iBakEJdFZr4nK7w5tVdojLZm9WGAM
rcL05Weq5gYObX3JorzXTh/6rmUviyPCrwrjvsA75YONVDPhjXbkPHOAGBABMeGy
r7X/Yy2RP3tG/DyY7nYgAWO38etlz7ppb3gFP45tGmQDEnqvttNQuvtBxqDFPlHw
gsDEuUNsHBZzMNgWy7vRKrAHL9uAaoZAzD2u2YZG4Wg1GWsn2HlxeRmnJyWDyHcS
UrhCZ+j1OrzIaLKgkebqPnurzfYVnRrOOGnpHiDrd/U5f2pDcpNvJdtyXoir8IXY
+LHY2uSOF+QYukfOy5WxY8kEYpiW+I2DSkD+e0d9BDYlrBhf9khC+njItJs8S9DX
UqpZ2cqKmH/udOAevM9azRmWtP/ct2PNWHDm6/nsm/sND1WkVmeYdTxMxLFQTZEM
nogzH3nFxflM4/2bvIs1lAwBSAHD76+vvHrZ85rk9w1F5Kv4X/HDLFF21TYc1udF
lP5z1pTpijQzk7/z727tiLajnTY0tt09H6UhmSKTpsugzRR8J2hCL0MP1PBTyX7a
IRLa8CLmk3d2815OiH3M2p9eoVbwl6Hir1+pffl5z+ROI4rcybseXXvlDXa95ZvI
hG4SwfxRlg3bRJMokE6tDOjBp2qZayYy405W/frC8mVHHcxQadqgaFq8prYkLkF7
bNXH0U4jX/ESV3IOerMlrpseeZ92vsKK/U4/OKFGzHdaokUU/HZJ+hRQN6uaRHk4
aEbyZidHoAJpDP+PJ/d/9pKBPWtRINIBIGMAviYsloIQYoWUUuYVjYddzQsVUlAv
vatTYKyuJiaI4mG4vhEmd46IhREYjU82vbJ0MrWds5iHozGTx03/DNvWRdzmFWi1
oJpsWqfbmcNgRRii9YeLcll9BCrbrp82+4tB+gB2tZlC3Uax/s+lUndvkrMejx9A
Nc+Kg+6418xZUxgoTrbfaLlfnVlQ6Z7jtwLWLA2QLV2DTOASQbD329hPweConIuQ
OMJiIux9R7WolbemAItLpjsB+CsyMJOW68tfRS3WP0boqhBqukkx7kikGjCejERJ
4oK+DC6l9luh95AIV7WWB1J3BVXMw2NNL5luCvhRzk4vDFytUj1aO6/yyRAi/Tmp
5qxWsvplixrC2sGvN3JvKFG+NsXaBZb860PA8xMTq52wGw0R0+ioJY/LcbHixcgt
kRuMENQsuWsS2W0SPkJDNRXfQsTw4Jz4g7BwDu7zjmlOeJktf4DRAoZzrKYYEgV/
TQGR8Wwp4oFOJCFX9SAAAw37qyvUKoYf+Gt2FBqPEIpPBQzjfqJweDvbZ4p62Db2
C5AH7AT6Joa+mYSaDvIcL+IzJDEBBSqk18Vb27wDxL/xB45ws64yNIo6ZKtZbxR0
gsMtTIj1L66Zf1iHJ/V9nzW8eW4qkYJMX+Dsdx3BNvQfFZaB7DKWjRE71/ajwzNu
Y4Duyiy6T/VIT7vf40kL4Q7HS2jwm0UNlqi6/FsGJG+V0bFwd8dlW+/ybRNImHSZ
HTAdSMsE8kqappluIKhCt1LNFhy9uBmZlFr1hI6BrqV1VnDQ4GF3u8wAzLJHV1/v
uebwXqGv/mSwHnlUppKoCPzGSTFKfzltxseof42vLrdBIFRAH3Bemdtgg6y58/fm
4OkqETvVrcTgdnVj44Ba2/TNuSLomz4ETnPTWFBXJmMmIjJ+FU7vi7OE8ZwRienT
z0pnstZJWUdWh5NeQOoq5KSQ6xZovv/EAg+80hH1fP9LTuOZxU628CoArk5NZL7+
6wbq6CF8VHkVEDK3P/s3tsUeXMSNuEUMw72dJ/gJQ7jxANr69EQuKVTJyh8KGz8a
kuCItwa8g/4qRWManc5p8Oca7dIVx/SeRwezCHWP//FQ4UAyuQYaKbx1x7F6HHhY
bIOmQHL1EAZSTfzKRDpdM5mtM6B22kBdE39lNPMp1l0T15BQcbcIIS6IQ3WWJI7V
x+UvRZpQR2HJ7LMrDBG33VxCRSapwg2zPymk6IGTjp+KcSuyGbDB69FJyNyclf8W
wrIQ1/wUdP55qjWJfhUm2L/opcWjcRvjlq2zQC3936jorchD34cjOol7caLSk846
4AZa+OPS+eryBhpoQiVezGWfs/0eI0okzPRFR7Y29Ld4nma7ZlFYM0T4bzdAx4Hc
gK24eFYF5zEVjQQIHKug+Mgh8umpo+0C99ohhFZHTZO6HhaLuTppb6NO35bCatm4
PCmAUN88uODVIc54B2fiTK2eAHQNt95/A5RIYud3phszbhUFLupFdLdFwsygvkTR
Rm03frUTVoXrmrspUQuSXx22KGmRe/WzNd9e0LHESwk+cgCS2HMNK9ceodQYr7NZ
9txP9r2OzwvC5mLO1QvXy486eKzJkwQ5cKAKEnRSlgLRIVnB6FYMEvfX3JzZmlau
MllXNU77rNu2KMHSun8YWs6+XXmpi3uXjbNSm8PituhI57w12f2SLOj/x+aJvVYY
z10YJleRJbbG61v5XvC613dod0BCFZZB0ZN/HG1mne8+5bDKlcp6yfMOdH6ay2Zq
I7n8kE6SaE47EgXQ96O/pMogcX/WCNpbrr78YLwHsAXgRlh0Y+I4UPlQmgTP4SIc
50fEaaBISXRVXnaYR1gGvdP5S9w6sj5nNHbkqmb0BO2WaRLtjhThvWE0GyWlT4E/
trQpf6IHda4bRYVbNYofoGAujtLSuExH5eILY7Jdu0aKeYbetEYLhJIzaE+oJ4XP
sf1Cftb70bTpn5DNEnO66023E3YhehVpQXBLXpa1LJNBcVbpgtYg52KDWzeolQzw
bly26qIGE8jixoC8L7AJZjA5dE/P1lPey92tMdZUQnLBYE9bx1IlINzXQY8Zr/5V
TgikRvitwfkToYzjQza5jW0HQY1XdPUAD4hYrFBSfulxvdd8X33eumaz+PfJlro1
Yup+HQTU5fzptGVsn71qn8ntcN07BVj7ZTOYolJ7D4xi96v5vHoZvyh0+D7sW7V9
VhXyISqTh4RQU6zWOWhKC/Emmr/Aw4Rbt8CtmZd5SxOFcSxqLdJxUXdvYgULzs6w
AXU+618M2IXm6pwGAVhf0R6y5ndWbh/o6+BvV+F6ZW8Dqs/M51f4oV8dDhb+DpKK
CrP0K7JEvQ/7AfBk+GafhAckUhavK0XHrT/ufc7ASFMQ/Q0eX1b4wrDLEubql7eb
pOSGdwKH9P9q3rBipD4A4tiDeAkq+bmWFF9/yalso6NuqC/XsSPs8lElBcLXltnA
1WtdGP0zSnJbOzlx3PYxVt32j9LcXNzPvffUMev4TaUTYDYyIKcWlucFryz4Fekg
nzcA65yQSvj1Skgk71ao74WSgzJosWTF0zxxYnklF3nuQgbs9nPejFl7XReMJbhy
pPyOCDUt9RKGdNxxPhfJQ0rUDny6Opu3qsaTNPpkTcxV7jdT8Lxgi6WMUfaQVGcI
ATGguCoq0+iiCuFIvzxPQQEyOIQfpCZCyzk/rVEinqID3v3WLw2G4qW0CaJsrQ3l
rbJoXmwmvkzWUEx6C9yHFcrTpTvRZikf8oLr00jMpPqarFayV8GyISIAYU2d1H10
H/8zEtPYm+Nxz/LiZMk1X2QFHpDU+M7F1DhRqurRTW+CnAhe/d9CrSyRxefu7A9T
MmYdeEICX1HoOGlx+7TacP4qanmSuz7cGHUdHCFNjH2AvHXE7hP+JnYBY2K9k06Z
orpES+od+Zht/jjVOB5mpOoPVHlXjhUjHIHzzl577FZzcbDcD1lOcazGQiH6VrdR
Dj1l3A+JrSK57WzEJh5bzYriJq2PyoGWjQoC3Vxp/rfUeEJsJAOj0hq5XyC7Fp1C
bbAxDXi7xUd9lnW/Axk//iz5bVpxPI71MXcloqmXQotQk/4Y3h86I1TbMWwGXIvB
zZbcRzcPppiT9vzr6KMgytib1u1qN2Dw/Np2fW6i5zzD5NFQCzvN4rfXBefTJQDX
Xrj9DupxNFJ93maZha/ExBo6gq/Lza2kySkfUJ68On68xqor6hpHJSC050UHAtK7
l8CHagCh08bm8dV8aJI48w7+91gT/NyU1tZH8kUWp3L1FmFwWunQbSXi5a5Wx7oG
hp4rmTg5uOjB1Ui+9ofgjdAP+npOs5Bz88rfk7N3vk8=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VYvsgmqFM0H46RnrVkSokhCM7RMc5WoQ+J1T6w0Q7qMO0q2wwQseTivUJ1dPcyTU
D2ZhMzCCsv6WdsqoYlCtDELuK2XFDfYvuHm1lQ5SAWVuKF0fsCXhdtH7UBb/TKVD
X1zDojBZ4J9sl2vF9mAF9CR5k7phel9p7UX6vcW1JfazMYYrtvorctwgScws7cXi
c8kz47yf1npO8mncQBgH+dSwhRBQ9ynkHf4YqLTXW9+qdNz/I/aRijhP5cMofoVj
vncnyYqILQH52U9u8R/jTfO3Gay0Vr/W6y7lD8Em5OBDjZxFe0VRiaWJM75Ilnwk
3BqS0lNwadPJtDItZXOlcw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 31328 )
`pragma protect data_block
ctHm3JQJI6qQCeqzMzWiyoNRnLEKMb5+kLzFcFSByJqRFUFSty8sS72zpv49i9eQ
LS83Ks3cSF7yga+vNoQRsYD4RTmt6/8KhQ5R7hyS1ZboJf2WEfCrzCc3T2vFq2gH
UAbO7O4CBKPML1SJn2IxRiqerbnuxc9WMnRnV0Mr3+GB25JbzJenz3PBQUeiMVBG
D/69e5NtIBtt+71dU6qT17xsOckQ1LiHIu9yscVslW9STgdy3MtfoioRN6XZwMPa
jDKKYMd3LU3Yc2NSIMhH2nbh8tVnVLdwWim37Eo/sJgkpBxzG833f+Lk8KhfByPi
TERHFHJ4L486o9roCPc5UWtTBOPdXSxywU/vheHqYYXB6s9Cqi/ggR9VH+xEiyIp
5OWbzSMP6Tge1FB+QOoyir34qvdn/GEeu/hbPP/7LpAuNC5oHfJxATcQb1V3Xhzx
vZKE7I0HnRb5FdilHRGq6Zt+7dvpqQ7KJkfCLEtjZnOnJrR9Vr2XwX67gDGmhlv+
JySJ+fkKVoiPyleap6iu5CAN0r7jUsSBphPYvtqTVIknOF+YB3q9B2QuQTzAZNAw
yjDqx3vwwT1vwTSIx+Sos+TgW02Qs10inxrLgZZ2ODqFJ+8Dzc+q9T/gqKUr1uJl
opsQ/3fFyaJZmNi+goRpfQHhhlM6J7UNQhHmQojY/6micEB13zTRE1Y2ha9LkHwm
hTpPlKWKWhS+1j6yiJLCoKzuuMPkems28D31eHXpC4vWznZDN1LbzR3dHmyBPTEW
qr/goGOHB8j8BXmvB01RdWO6b18yo1uHmL1RsTolPAO+8i88Uja6h0DzWop01Q6D
pnkMGpFWD/DTnq60C3nYM0BG7M3QDI6dWjsqzzTmVq9n3UyQtBf8DQWKKr/Go8/q
l+VqlnIj0tcxlOJh8D2dm0kpGPHZD1Je3fFRBjAkx25hoIwN0nIk5bX2YCmm4oTA
3nSmBLARBWk0vSTFuNfs3wIqH146Z/8lAxdps7OeukqXxXYwaBkyZEBw0pXKAEM6
IxwERVsEpBAwgStXaUkg5dleAIHrhYZVSMopUlGT/ziKvDZ87SS97lH65a7RP5bX
TMr8MNChrBFvQMIqhz8l7e04HCJZMbR6slGcTNu8nhR5XwsIDdZq8F4NcxYYxB8T
2lsU7+Dx4GBLD+ALHbDFcJLaSFbTyOAqRv/nebmgBQuwbHyNsLe6SXZ9mH0YWw01
lZRE7rBTis2oCOk6SUXmpQyKAdfkyfHEZtTD+MIqjKWo1r3e/6lqGVu5owehsR8c
o7GWtgW97E9tDCVkjq3JMBWs08DGKNtC4yJV0GjHdrY73GiH44YEEofa6Hk8aLLX
cyogBFUYDJTda2Ci8wcxZpCqMxaQiEdtCr66fEfdHv33PrMp4SW/A1k3u3SLr6Ze
3CKx5AIu8Q8om2LhnaOPHjsVr61Zwh2+Sx0W79JDRmOoHwN6iwLQsw+1D3RVbiVT
cGaGh2J/2iCLR00dF5J1AD8uFnskJvldWrwQzBEgNvfiZ2yX+MNSmonHsT3j1tlX
AQm/oxkC+I7WO9lji64vh2Wt3tt+TKkVaEJ2SDLJo4CJpRFgr3nmSXE/cY25vq0w
HkZVcU5ifdQxN1seEzHtd73HrDKhJCCpfA8k+oQ/Lnlkyag8P2HRH6WqmsyqDWRM
3JencGLSPmUHUGUHCOIJnTbUNsEOU1HOzK3/uxfk+J2TeBCJjcwYn8QOENCkAEkJ
EL58CSxdaZaLLtXQ2bREwPYZ3Ism0r/it+y1UWLJh50SFwGnzM0mY++wDS3o+LRD
gojG6WBy3xBnb94yGAG33uttOQUre6+u23WHIt1RgkNbdaG3rk2vGGuFFW0TVdCA
oAU+jk37xi5jkZOYHeG4BAaGXIfe/E3v3gA/wCIB3c5dqeh8jQG92QvH0WDba0Tk
P3204W3sfSvJBcZ8Tlj4FhTzOThezumb5RZpcyW22mSX7nVFLzAaKFLo/YAi2NkZ
LkNg7ZZlfpw3hfmvwUGlrOi+xCzGxecfWZ8OC8hj2/zSsWkOaA0civIQ4X40Rfxm
zYsrRItm5s2P0pxr8YJVOYtihzYP6LY7wO06yA4SkL7pvWsc1HU9L3/xJFPQWa3m
Zws+DXEzLtn9lvdt2yImPqfNPuQTAmW+x4luDCyjtmiDBR0gKH9zZCQ3G4bcyi50
ui866VQBLWbcNYlJZ8fhL/L/6WoTfpcC2F40HNpLE0nssUT52jIilRk0iznrEJmL
iLIc/vYJiQUsdb+FCSZPCPD8PSAdi7nOsumThFHA2p6CCJkCm3KkDktj8SvTX4qd
OIMeGtWXUR1eakEM9ifu/MWaKIDja5AJjXjkwrxG91HBihbFWgqNn4bc8K4yPGST
5XnqIcJmaDIMPToCfDDCCowB7nIP2O5JxbZxlVu+0FXCyray1tONiaEDHL/eKQy+
8gNgpFRrda/xkb3HEOwZ7lyHf5ct4wcjmRqrNOGMaIKBTr4jqbiFL6iGMiP21EDO
Yh1nlZ5yzb4iXbk2cOsZk4s3x8cnJ9WM2Twn8PrDYwlt/4V6Y7Euc3EUQAsrylQ1
x9BnRAIoxSRFEww1HeeDCT/USDWDl93mWDSSdVUICAGy1xCrUXyQ1/X01WMBLF9q
DIiqk+/P1oVTGJwtny2uqHBTWW9Rfi7KdALPruEx+uz37RrZ+84MKpgiC9iVomIc
mPc5mctOp+Po5N94lWtU/k9yfUyK2JFuQWO2L3BoZw5naWOHCxQmFa6vhJta5YKl
3TPU4gupYimTtQsC3HG84eS3ohnIL6x4HtclX5LHRZwvMb0SgsgB7hKeRIUZowE3
9EBo5X+WQm65zQ6S7wrcadTNOqy79lUy2FshmYPzZGedtunuDysIvtZsZFmbp9IM
mFV9DLzeJ6oYpHH+kUgGa8CqewDRONzkMl8xi8r1XwTZJ8VqeltyLsvL1/0t4TQr
uyUAkzJfaewsq3oeyjittFhhWgYtA11EMfukVh8GLZb51lbFaWIiv87iM3KIIVC+
ek3/G3k3L8L0NY7X1PxQ7P5FXrsCwvsfOtV1kzOcgLIfIlpwSQQZz7ASylxYPdaG
mCYK6JEQyTg2y33dGXjlGSUFZmaJj1RqUe9Sk+NkZOBT7F/WlkJD3NpA3VB+jK2w
DwVtaIfgbdy668ipZ9JahZC58ob9hPgLN4vVJe+QDpkOgXR3i8qrEKrkiMsI+KGB
b3ux8/FOf5C2v4Dlvsx/y0BhMMIciluNbzkex349EEvepIJd1A2m5IVQ2Ho7ciYm
VsR+mVvV+9F04MlfocHZLUjO5b/wOz3b/pAbrlHJRHEoSSmeGId/+ahU3rI+qv5d
oMopEDWYrCHdpOIMdz2PfnWik6FBuefbf0JpsJ5Vu0VkGD4vaTutHCZ2ij3hHBi3
m97FXXh3htXoYQzDAGlunaBJ3dNUaDl4OO/2RkJQwd6b3uQHiRbQMPXqVx2BF7t9
grQwDjPreyTFdvr3bjwQXjL3aOjXYfup2WqWGSfB3Ov3RZ4CRIRQgZA/8IToV7rR
kt+3yFfyjpbWL8U0l8jpzos5ZRzLmbl75ECYRuA60d1/pUXTCTmBngttAYN9zMfS
CE7JnE0YEvMTJxpKvKDWZFWLC6xOZsiSQudGI5fgkzIlZ8YKVZ8GX0TWqsKWhCP9
l3hTxWiDBuWWsAc+m09fJ3i4cSrZpqNlEFh7qJsL5RI/ZHUA3qRk5lHKgf9x2DiT
ElEnTbDhSAyf+WbMCRwI72VkB74mmJNJa1x3YSPmAUKfIY/rh+w6YBFNVqCjpbud
+JGPikqSJmOxag+qcv6mgWRlHzvVwzu/dCuJRhljYzhpDxj/6WoGk/gUyDwBoU5u
TlGT4aYiv4HkuUw08HK0rDIVlNcz5kJFatU6/UXXYPHyl7ioK6rx2Hl/YBleIUGV
Ydb9cQBtRMEh3WWbB3nKtxUPuB7UDQ6rfTl/a/J7CxledPyCmSEPX/sKZ9Gk2lsq
cKOZJC8GXpzc6rMT8IcOUn6kuuovM6EqYAYrb9CZ53+WNvLqM5zH7melX8BREHbR
on2Jj2Xe995d4Ri4+mUsSa0nMT66DvdrhDmONTRo86Aoyu8SlUJpV4Ey2vG0aLRJ
qJ2WQk0VV0SsNEQ1+Vp1kbuH+H0qg1pWO62VmIcrZVXQJLuL7NE3fbHi2VHgGRoK
kOGFbK1+6Yf/Vasj5slqNv4FH/LPeYjB4I524NcdqFwFImcpO/vOpeBXzv/myERL
syv33dGpBReBBxcPO8aX/899y9/NGw+qDVCcSyJx3RHgUY8Gbli/2XOty73hpNxL
qkTLBVMJUmLDbzZ4OZvOBTJVj4UGxQc452XcutyWnCxM+m88w2TzOaSLvnnKAzmH
EP5TxD0utGg2wnki0XEzDQhZJcj5KobsJkWs+fa1EnvlebZifA5n1dYOd8x1JT8E
QhG7PEv/1RAM8elfdo3swUFgFpfPG6mkcXeoRk0NWjJlh4XHd3iK1XWiHcbSyZyg
VOBuNBecek9tMQitZSNUWuAVhAZSCuBzP3EFc2zi8P8T5MGAd4tEfdeuErYoRN04
gJlN9mGmCH1eZGoWnYeRDdmCyMSo0pC6NEbhA7ct//NODapQ4RB+ZWcuG4TqV3m+
bo2/kmpj/58yW9ODnvm8SVYt7tvlLJxASWTLNggvKXLUzBRB0ZpU2iuiX71q3ISI
xcVBxS/dnUSo03vyJ0DuvEwjiOjtMDG9DXFhDcHJGn+HFJPuWeSKSaBiSaYZ2o1s
3GruEtUsWzkYHg3p3XBy6my94AStC5ZLlQdFebBlp9+piWA0AOrNxU2Z1oIQqNsQ
OWYI4MFkNvJUT8KXsG16IATZ41+/V2GZe5WMzLnWiPs3ON+jUx7Eg4eIpu4PtGTt
shWJXQHZiJNaz6hLAC+zqkjP0s7q6Dc0a6CFoyO0akkSJHr/4z+CU/PXF3JUe47d
/kNGLca9qmUrQpkUKBdPBLWxAgheeBNwKUaD2Ud0z9YqzxW/lFKUOxFsfhSvOyTC
muHcWFz0/OzpiMC5W4eNBRHSZU23StSFGi4Fl+eAimNSlYkgQJSCTIt0CpXEEqXg
W8OGflX8/28ZTwysQszWl4SinUh1UOFm55MLalrj5RBtzf/ui83TM6oi00xrhxFd
9WD65TQgrnIREBYiAyLscgCIR1UZoHwxoRpQ7CYvd3TbOSm9GQI5KD9ULOajW7/j
v9KQmwyoi9B12XGCk5FzpuGHbLRbEe59WlFF9wRgEzgVp761wH6CCJreaU4dqW7D
ZeB/mAkrVYSFuZ8HHOatmeFEkw4+uhOcwBdDiN9+bC/zNtSqkL+IiSc53rkk/gsv
3Ho7v6nWYLnOn5dpSOlPcT17U7QPikONVMs37Jni75ZYMc1BsEygs9fOW/Pl9AVJ
TW061stRw2SP4s3Lw5rlA8NOtcF7P9RhRD2EbyZWCXpOd1qYBNvraWZmEAfrrcnS
CbQeMqo3jV9YGwZQcLFCmySre/XC4+u4QDEOue4f8w7CMlj2FT91tnkkve0xYk8C
ltQrOyahMEEhjqUREtp2JnFSjY/Qxj0HAaNpylrB2PCfZEfduhLi1/EnYdoGfjJm
GLoWgqBLZEKocf6TTl3p/6o7N2CHEvikUrFnbJmLd7n2yp7RjmILCXMbXpl7YEMO
k2Lwfnt5TACp/phcY3eCQhW1xjZEfLaK/cCvi0Brnsa3pGORabkQlAaqudND87tS
RXZgWENfWF6fjl2ArDrvc4sT9MPbMNMYfDe7Ub4D+J9ImHOrBtEY2podON46UiBy
dAjr6f/thmYjfpE1jtcvPA78C00oZX9OLm8AeiSWXuP8twtl+zOpzxBoikih7rvc
BAt2tWG0odrQFsFK94wlanqWFZuHio2Yl4dGXJFMMu3Vatdrolo9QkRPTBuYUS7e
TS67trs4E83NIo7i0s/X4mk8aCJSGEGjGbOx76EPiezpkIYBc08aG2S3jZ29lUHu
yq/HOrn2el/YoKhaMrv2LU1Fe4/gqh6xqbvFrq2jV51hBOgo4UJeYWUL9EPVud7R
eKxh/6yFdeJlA81E5hW0FanhwaeRo3Ya8pamKi4JPjhXigCIN4x++1YZhfyxoMib
yE9WOXUSxBRvEMrsySnJqnFndcjPFPU/dXJnvQaIdxqmSqW7SBTNQnsGno7Uhkrm
ZSimzOKiWWvJkeKRtRvBBIW3TXV7vw0jbjHclCG7GfocwTFbOS7ZSzuETjRcQ/D8
/dZzHuoQU9CB8pZ1TYYnw4vWj37qq4W3DEGChU9GhEz0sO50ctuOd+hrMn1ayib2
lnzMXH1mzU8xjJllMt6MV1OqvrBKjGVD38mp0aofCGyS5P05W2Al1SANREXoKNNH
r7zp8dQu88nzJDQdyI/GslTdzM1s4VeQHGiyzJg5vafGnhPbaWIzmiabirw//XfQ
tbm1LtXGuBH9AWuJr6IlqnoGR0CysBMY136bGYK9NXy713iQY5e2da/baBTSgk5d
dDplXEW+wVlZDEvKRkwYoMztSjwv0woy8cF/hcJuRepUbAjI90pnWMjw4oH3L9GF
4oKlZBYRq86L1CDbT51RcFE3HvQrvV5tpoObmHov+OZl+Dk7xmh0TPvrasdN8Cnt
CVwodmKHTD8DkFrnAL79kn6NJoeGGzS11t3WcDAlxrUSdsfOzIHV4R5z2ztyyp2a
TwM3juj66BvIvhEejJ5hKiudsnTD2Mp33Vjow2BuqZF0ZdkRn1gU+bhXf0w5KD8O
BEuW0WxbWWIa/rVA0jXprcuoJU/EWxcyiAhUYeWp+Ulvr/5E99u4jVixXUIO5aVC
cth/eqKr+G9VlOpaU3ky2f1lQzqXeWC0HHuEV+vA8LMoMvMlazhnJ9ozF5DwzE7N
MLcHahdDN2CSZwSaVEWcoHI6ij/QMpXp4zK9byhWsVnMSYChpGDBGNUyXKS/CneT
4H4TnEm5Ux9ut7EjVjP2emPsRci19/yiuQhxw8qkpIS2AP6FdlV3fmluLlIh2o3Q
EcsxsxOaxVodXFNdmXlGdcrRe7csPX2d++f+61Fz3YWRC5dwVzywrVxUFlXFu3E6
5OnpqBhOlsztyhlT1FK5cV21BxCUvhqV/oAueuGiGT2djonwa63icOEmjZIIPKbO
JWQ7VeXQ7CBYYrf8IepsA7y6zkQWeUW0/4CbVbwzlpq9hMAEZ4bWUK5RWf3agc70
M9dNr4sRQuM54mtwU0cwAWj5DycT+BXdv4MrjtqPsWZ/esVoRP6vhJv4c5er9ThN
yAcM7E2G11Ak1/c6W9GUM4VJIjR9E8OnwRmH2uThndOgN6TBGj9AedDEyaW9c4Sv
YV3XCRu+M4c18F8a5J0qleyiPZujveBX51Zld5/5+sLujFnJjJWcbJpD/TfckmJu
UGQCu823Vyc1GG+pwGmdgpWkuxJsExdf0C/D0ffHaJca2jFQ7fQnIgFawcylrV7J
mytLFCm8xzuLZ4spkST/tVFvcIjq6uCkw2VyttM/ryYJHOA0sBKKO8yQmOUwVoa0
OhRq+EkybUXwzlhiQtZnzzfJJbObcM4U9EhLcksvziRNQunu/MydCER0BLVFypOM
4YCW6GablQAG4NB1errhD5+ZLVUJQNmJ8LLRdjR+0YszhSTjy7RzV36mt98PINyx
M0IUD1e7w9mklKS117FAy1dsHrSYB7qiT4jhNGtBy+xh3pbDbgMpa9XAPXtnOKe6
cAuG2JyO1fqsaeWIf7JdwLMT1zL6GI1NIT5IaCSHloHOpgLAdFmSrZx+uXVgFEbY
uG92av913AzMt5wW3/a0qfBegPEKPnJPW0rhHqqw+j9U8CFJ9f2fQdtrmzPWpVe1
3BlbGwHM5ArOETsrQVJ4U+J7OK/nuZcIRcLgKEeqhO2E5kXxsiDzB8j07+cjDUKg
ygCrDFhsbscUmSpiofScfmEYkGMwwNNesiOp8+oLHH4LO6bTht+iTHgtgD/i7Suz
7eCAonLwoufPqNdCvFeTBDpFf5Unfqlev2CY352m3AFzDKksJEv7K09D0AUJLxFq
o+NN+ga0U9VTw8wgPmLExA0li2Mh5LgtoqmGrAuiRyFw6BQ6p3LJX/MN1X84aLGd
51xVqbRVHwEVoKWsN716620wgGYRr1GwiBu9XRKHIO39po9I62LOc15VPY8M0YYg
mas8bpUXMF3ns9KyxhSDOoYOo9T36s8gfZR5hiIt7T+mYy1E3VaeYQulZtUc2Do2
MH6LVurDFJxUL4tluwCQxxckh7MjavFVSTiz1ma4VSLZ/89fhtbLHdX4SHtuBMCx
+mmzMno4iHp7oB5pUqVTClQGOMzOppc8G9xrfMXUA+xdBY7TBccQSahSPfhapPkD
Pcm43EPfj5wVzvzLM6AyoJSIet7ZfhNtrtJBBbQgavnGtZl/GXV9a63BYzQTIRd/
ImWy0GRP0+BzyoalMqdDLFHS3WN5E3bl14EOfI+KR8dKRAQiLNKcla7D6ShT1rag
Sbg2IUw2AE42IapaE/AKjowxPZ7l6h2g4vIq7oDfDOrbQqS7NoHqU1iQ5QUQmcf9
6x3iEHehJn4zhXbm1QXMrFtRjGJwu2/SUb8ukk4kYnIodJIYJTZIR0Oh0iCFTZ/r
UMKjOTZlAFMpy0eHIrzWIKkHzP3x7bDGs/hZ04FMBWwWsD2axiEaqW3/0O1jPB+p
CDlUWV2vr883rBjQSlF6yd2VXguCyMU8t4kswCrfAIP935qXP321ByTZimGpcO20
+lzfTMWdUxHfkDnbdHryAN2aoPmTm/LgyyaPTwm5BfPC9N0elVXMq/oeEcXpBpVR
PS9HDLladBQsv1dKjwlmPOkHxEL8uvxCGSR5Ub1Dj8avYM/SxVTu00CfhgZmnfbB
MK8ZcKnFOpww6NZVRkP+JcGRLwq85lwvEJND+06yyrMjlZJq1CShxJtIrFLbtse5
ugUEkXx/fYUQ78uD4wW3ZwUlWbums+Yabz+lUHcJbB7746UH09q4xAh/LfezV+++
VZzxekzUqseFzNzNg1rLctrVZeKCwF2NhTdFotLwz/er6FQr2IQNUrn92GLf6ekf
Bl30C2TqauaRt3Hkj+EceemidIZNZFLxXrUqaJlquZve2IWSZmLZxhmniBbzI+S5
1ORlfPjzMsurOKjKoFT+1NBIULCCMVtYOnk7YOu3e1B1bqb/73p2du8pxiX0sSEu
9sGNe5qLcFrmPvZni5DDmNontf5VFdQ84QSSbLzu3rDz5JWLsvc6mqVbdJNtldiL
SCw95KQnRaV9y3dBAscgWD4Ol67GlH6PA98APT6LDayAwR5u6R4nK8RPsMp/QCBn
XU2w7iFleaWkMnJK5y8I9LvZoSq2xDMPFbe3JKIcyh26GMxXn6a3iw7Xp+2KKTXf
b9hbpCoc/bKvAyza7NvkRSJM+MXR98zVTLOOk7m0bzlNyqlVHrGz7eDPgX60BmVH
JRZvAqvjkDTQT6zfxfP0C8skLr7/tZahrftghwZ4Rmwsqf25ZFdVH5ZCA5//ymDE
Y3VhS6hll2KYZLFikOFUrcoUKjaoccU5lUjk3Canmuq5nG4EpDyp5Z7rHD0C4Mfo
fa9mwf39v9plzPR3GFPV7vD6KcEfnEHYJtm7X/0TqASeKRYT7ic1Z5ENdTTA5CXl
V6g+ry5a/1qozS3bSQe23qKLJaQb2oJdOLs5HHvQJmJyN7eb/KTqRsUZC82dGF9c
L73UboKnMcs2H7+NsDo74Iw7IHzar33aOnVxaOFe9kB+GhAT2xQOTQ+G7RSnVsPf
aShgzY6z3d02uKx6iP4MlxYZyxk5BVB7TVKtuE65NIf/SPBCMWdXS8DJyr+zSEK2
ckA7UuCavKWtGhTb+5qZiNbqtog/ifR+z9fDe1+ZoxSrRaLZuEWzxCruIbBpOZyZ
M243fqZ8Uj+nLs1ATe5UUXOeEcjFtU8CLAd82WJQxbF6V9bmBTadx95gzR/lfWJP
dhYCP9Q2T87Rgrbu8d6qHe4yoGc2w806tZbVdjqn7pK68TgtcbivpP91//5nHrfg
BQ0AqXbfJEPHSAjeZMWwH052Cnj/FoJ/zSB/Ww9b3/qnq/l1lXCKW4D9TK8eOkgt
bpaPLZ+/zWTjAeod2YlrMfGgM+2kFntypBPbV5eH+jAnmtQm15J8Oxw79V7xQEbt
mhM2e5PjJ/k3hmzzGi21AqC1fe5004Bi1jchbZD/SvehX5rWk9txgaQeGzQCdCan
RGjrQJxPP/UUrMxtpkI3xOKCSLI3y+qC9uHad+jnWf5UEkYy5r2pLLiVxvOpDHFL
EBQIih/dZL6zGVa6biqh1wQ2uPiNFLlWRd+/rB3c9FZAgYQ0e/wAlLKlbtUW1eRQ
4Eqat4IAzjt4rJMRANgaCxkUcEAAuQyT077DwcM4vEBxVHOiYxDqqXENdC4WpzPx
J3xv9iHEUsgpzlYYS00kf1Jo6HSOJfFHGD6ILF9H4qWlNGVeJA/xb3aEhG+0zFZE
tmWbN2ZgIwEuZyFzhjy/CQ6ZlxQy1Ki7MEfhVqdLyDsgiM2HMr/2tLc93YlHxphq
qgybZYF8GL4AhYD/UNJsPwsCar0lUjnBeps4VVX9kvPUQSVy/Z/CoC1cY/jnD95I
+W9+yFiHitt59+b7iSOAG9Hmiq0QyXMkwzgpoVVSXHMxiJxGyI1B5CEMb9NXSwpr
xxuE5dsRKesQ0AmzIa/Q8gP/b4hz++ihPxXS65P34s/X03Ee++QDwOawDTe2+MAb
PiIYKJZ3dJtVgRHmMmMQrkuRdE6/YY5WMo2/HTmZS+c2mKH+/Ew5qiXG9z2HefgB
a5flcxSDElCb8uL7yOvk5jiJSLPG+PL1YgIYmh0uVtxvf8YQIFrUTH1Sg16kcd7U
CRBXwPjG6PpMre+ULSWYdaea4iZFL/OMBD/xqft9sSuVY6kpzMKIVPird8vCOo5z
fgqX9fX/B1goDUOaDsh61gSzJ2JwKo01hrTrdiED32JOZRrHAUrygEnS/EcYuzjX
HKkV4KtEoV7uamnprLCS2YGVfPTYRZ0dNfRQoVZbSO+9gRcwr8M24ZCO+FKnSbuQ
/j4GO0KpPLYku/VOW1VolVaeoSwa5I2sNF/+SvY1AzGjSiIVvF/qjGyehPWDsbGh
hsx6E3fM9EBKxHxTDijUrY4uXHf/1qABWhxZBeYOh1i1QZUvg5xrc+IGAG/xVG3R
SV9mDc4fxPkzyf392tmhRnPOJ2kbAEoGK4041Y/Beil7JCnQjkogrJanstlCl+wi
YMoxPcpH1CMEY0MthJVuieUYbty+q0VDyT7+l2w+z1xrTwtU2X4gxsbFZo+uEXEV
4YXRlwOs6sMlcFctwiti+fdj7iaKljCuNDK5WCUa7KSUCZ656o8Onwqreho5yHiU
oSd3hmcd4FbubGcwkbyhQxsQ4rjud2qA5Xu5poiL/yVk52wVTMD5aIWtEn4ijZOg
C8N6V8+tvgnf1CIR+HU4pP3Zw5AQwwIyiLMCkR2H5fHLaVnR/2GBsaJviZ2ou6pF
ZwepGvDcHmbms9HtxB0wY2IvPjl2BsA/0vLsJm81pKI1ZU3RPva+ztlA5t7kiz9M
Mx8SCf5GCyu92eS87m8D2UdjikfcwGKYb4MPI4Mw44Qto76ml517jqgRI6O7HCFs
E5T+rK1ih4FUKPF8/IUJDasBZ5j2UfB7qDod0NgWCC8OSITawTyEwFXHL3+vwmj1
u/RaLrPfPvUyJS2flFQYqDi10lD7C8Og9QEeN/0O3q6YbeQabtLOJKKpYDfb/1dD
SUz+DD8NvZvZaI4/LyxS27lOdoaFCXc0UX7dywDNc6g7UN5GOZQtLwhkgNgKKYjm
BLvqVpNJr74YzdXtQNMZz8Qu9SFn14q6SfHzInsmPZv0AsgOzxKAPsudKTSc9ape
sFtNj0A5Px6jqFIPwCeHeVFHxW5xEeuD56wByavWM5EDBF9k5NWQN1jJwlT5cSdl
epCIxN9dt0YnQEI4xQfqz+JQAk4tUGh9aqcvMWryQBF3S41TWeYBrkQzDyaMJ8Hl
L3zMzr9qvA3LWhqQmtvQgzkFsHJkuRBkwJ4oGmxo1yyPTW3PeYXi90H2143T4hXN
eDPeRoI758qQnhtCCI5ceMcfSA8pgORkSM9cBLCJA8RFTAixnCMKFC62bAZvj6hc
9MGi5l0HuY8TRmgkhtJVZyI7LkDJsFzo6+Wmss9wiSIb2F/O+P+h+YeY2lF2q1Pi
ojDAyRlMYqCqQhFXaawKP2PxxIoc8jbtnWCeoDyfVNM3jk9wQ6/wOA8M/uBt/RnJ
06Bvr8cgUntzA1sLqqQX9OJQKtR0B5A1+74kd9mgep80Cn/sGCatyG6qmo+ttYsD
BPel4yX2ScvlvbzYL3VVd6Hxycu3sTyJlkwSanDfvvhifIFn5ODzUNZs21Ehqp9L
xFPKU8zYriG1KCvVmpmk+Lq6s9sp9+j7+pnZIRn+9rE9NCEtnZZ7UTFZ2UR7kAfS
IFkfd76rXevIX68HTbiLEDwPaQHvLlVHjJJMCOGnArMaJD3pz0iH5jWf2dU0SyVf
UcTHVbS3iTBNBzrXcwZZJyN5ieDF6KAmaYEzWUN76OOY3SxNR5lN8Qog6qRVvQ9U
6ZFSqbOY7OlMoKcqa9sv1CJif8a/rlb9ashk+6NJiW3LqQiKpmppQMerl5fc4UhG
FUMf7WQyIwT9ESFHth23N5bux2VzQTfBqpqTnO/7Xrs11tAgRxpEP/rMCEqj8CJ3
wnLa5nbxWNF2gpzUy0qF+DsEiOFHmRbVpRL6JTDKVniyiSvt8QEbAypZaTvMnO1Q
MU4O9IE6tCtd3YlyQ8qcT1A8oLMeqK+9YyQp4YPKB8yZ3ia8dAofTgSfT3zTwtVE
K/y4+F8IC0Ondc2wzB06eX9o67eVIXM5D5Exps8le9j8t+jv+3Wiui4H2Zxt9IOm
nfxEfb1iAx00Nw8eW/n41N+5sTI0rTRxfdrt1w27Akahsqr2MSJpB9VO2ERzo1hk
rLU+p8xpNulDAUagJo8RHCNxHmxIpWD04B3QDzYbX5FzPPdRxVfN2X5Idt1i3Mc/
Rah4FmD6D7lCIYWzUuSK3xf18f048d1LvuxFc6I/87WF4awB4MeA5d2qO63ZAQWu
N9bDSqeeThjMICxUdxZfyE2NvNd34x1aoYdJj3AKVpKXTk7Hd78t1wEKBQUnFC+y
iLl8JOgcmafb8cWJfcz4i9sxU6/gH9qY2J/5fadjo5FEsp8UyM1k9IdM1rfypH5c
9s/kYMODJGOGqpDmEVpIrbj/kiL91lxsAadetGTxHuvmNNkgSIDMsTvybZvJp94M
R7xK99kJf3n1Dq0h8EIs37v1uRvmHcrUfwiw//y5pfi6XfXl/2cx97gRbIMYqVUR
2a73xdXTb2grjubU3JoSxDTiI3NiVlI7hbryZ3gDejsZt40EMDpFd2ReH919JUPV
9J5CZG2lmaFoh07u7DTKZtLykUuu1DWtqerKkzPtostsmc3N8kKjkh/1cidBq7vR
OTG+4TSJMQyQIFkcSAIPiKr281nX7S8cgA6kAeSmUm1/+IuHdM24VkNnUP6f/8z+
S/AwI+a9pY8+BsdtGaCzKijA4BOmpjpHRI6xiLIqiUaFBC8nCEwSK/s6chy9PJJ8
m7URCXBW/yxXqdlvtpgcxbMccIx6a9uGVoSveLLYAXlUnZTGOgXKSem2VU2nb9P9
YmbzltdAJrHTwgQh2cb7VGQLkiasrm5WLBgMj+dPwCzk1UDGbEPwG1fh1ZGeWulF
839xDp91y7/0Gqawd6JAFGcChizaI8eOwABLYFlJYS34PzDEEFvEqoHOddMmgxKM
uXsw7m5cgnlk1/rSJLxhnIv6dRsQeLipdJVHNqwKKtr1FsF7l/ZuniMidozgXPjn
zeqdAPzID2aZTwBdbUVLOr891eyiUN1ca2i7VPKakKaEZi5MmPreCWOuUETJSvBM
6HZ1rbaD+7KW32mKjewZ41Y1ZhsWTFBkPRrJjmkAVZpcQaBYKC3FiaTsrUXYnCEO
we9GfYhW9DjmCe1Xf/Nh2hN2Ju8Og5T2RvbKSlnAjdw8FjqhUlEn1ZQ/hI5JPmDX
Ujdy+p6U6nYXDHMvQkjuq1ZQmU8/h4I1VlaEmpTQ+2/NqTF8w/az0hFTGb0UbyIp
gNg3eXHsE2VEfRx3g+t0xZYWOpZB2rXZuJUg75gl0UzHc1DPu6RgAzfAs+8P2awC
rOWRSyISpo7+EM7/Ca8yk9mbZYNHctL7ID47WYJ3jNYE+tvAXMRVl9tC24uVU3Vx
0AJf4Dd4q6Et43lyYOVI7MayAI0RwtUw76G+b5nhoaKO9NYmkOGG7ejHoBxs9gGG
SdCp+JBCascBTJVBGqutgti+QndSFJAJLfBI4j11HtBaBHz0b+tOnaz0jq11JPzT
Szm4R8euoI4I67NsG7RSohJXsZPNHoSZMChi/GPAJtye2PqcaqE4TjMukDJYlD09
OpbiYeaUmG+fmFSq/WxDc+bfiqNLNN41nIW4G4iI0XdfGPe4TB91PyEue+d52UUq
Ce4nq9QmE4POf45FG8WfYMLAdH3ixSgfpsNEDKEu+TMxo/Xm3WyhsLaWGfb8u4xP
oBf/S3IU4hs1mlkKK7QDPpNHEd9BCxzpvYS6ujQyQqdTjdRtnZncCgVcfedx5f3F
kjkTe+R1DQb8x6wGgNC9Bf6623CYAHxDcrH0Gm4hzGRCyHyriOo9YByHekTFx5U1
Kp08wnsUVZkSAdNOBe/exohS3U5wK6YhmnHfAPdirc22JzfYQ8miViAb57EN+FIv
EJu9uMvDWERhweLMeGZzOJbCMdeysNkEgNc1OUL5e2OT0XirW38COAhYDEbVG1eF
qDLucvaL6/Gm92EA0jumiCfCBljC1tvlUoCr2Yn2sN0gOsYhUI9Nu945VVE4/3s4
qVv/hMKGWHwhiRjxnLZo+8iLlc6F1JuIjcgTDE6uO/JudehNjWY6QcZaptphPZxz
fL4y355ujH2kTfxKkyOaSopeNMqieReqHcerujQjJCvAyEWkTadu52aLaP0Q5hhC
HCZrfzxsR3/v7FRbNGkGl7NL+0Vwi1Ua7o0XqMsXghV1X3hURxfp9wQwvjEHUqB6
cb6ivoJmrJ825MEsOpeDoZ9KkctTTJVLrVWHNoyGbaxks6athq5WozclWvFEIneH
LIk3N4eniV/F2/FDi2ZZTs6+D9XD8BD3rWju4yzfVIvEgRNzCGsLxhRFbwbWrok2
ORElrOQnNus9K+AlLL+4WOYmfje2og6FXnhG2tVDbM6Y1oiQW6sY7N5Cja0jSDlY
aAdPVIh6fxPLyQP9nkWUAOdVNQ/I/yBivLKoUau/LOeGkxc29OQ1TLP1GLvcRhyq
nCqGD85hkQz6sooMCZ6tocScw6yK6rMBPk1KlPjHJYJ0Whe9qckPAC1HErfM3Tgh
HcMW5f/51a66peaTzBe3ki8WIRekurbzlkRj4q0+45LIzl5k73iPk2zr3p3FWRWj
wEPNJHKVN8bH+ITm9diN8zahNk6Z00x7i18z8PDbCsYaHS/6NYcgl2efK5++UwRl
5CD910KDL4XnUTCvMaS8GjYRAOYDbfG+IflzDqpWy95EE+0PJAhVtDluMgrlU9F1
c5ZKfY9dXfGtVSwhy2kcUFMa2qYjrZ1Eg4ECNlC9PZXdHxsu7nQ5YcVgM/5nPYJS
Dg54eOz3lW+7Cj29R4qVh/Lxwyn3ZYd2BeYvIA2+j7YEBA6Tvjsw938sNr8kV1zy
LKJ+9x3U4F8Xsm+RMyhBAmnAxfBofkm4OjJpUKk9wHWqZ0kUWVdPziGEeJNtgtgS
k41jKv5SSYCyYE+t8kIL0u0hd7TyB7yzhn5FeviD44O08iPdHcywVjN9TKNWMy+i
MVfdvbi74h+JzvWM/8JfaxzintvvsLHKoTynX5TjmTnsqCE6r9wsK3UlEjvfUcis
lnZAvn8BYJWUzsWPr1MozR6/tZep4LWtNrB+zlMMwuF+p2b1Gb0zGA+gMgLJcTk9
RLbTZF085EIQ3OFz6ZA/WrmnYVH3NiU1csyFFE8fR5MoG2BJZPMb4yuVkjxSBsNk
KIPuPTPuzOPGsNOeAl8kDJkJA4BT/H8IdZGmSZhLwgHW4DmLC9Qf/FtIdByLjle+
Wb1t6iN+GhLPbPZOzQQyMDK1YWghhO9IfuT+wuIDitadOOdNS9/bshm8V9XmxL2e
EpCVt8nzVrj61D9jg39DsB1ihoVlJbpot5EQRTioyLTps0izD+xhfZoDK0IQr1TS
gabqMh0nB00abm3ANtCcCVUcHpM2eHtU398cUUgvukCG9x/vgrssYt4/3X+3FP8r
P/TRhW+yQaYVnreWlO8G7Y0nBIDTIldBjPIpzNGiq32j/bBKGXQ+kx1vGGetY5vZ
UT0m/Yx6L8sgQK4pN5oh3YCYGdEFSdRlR6pYSI49Vout+PBBsLDjPgBzCOsCdwMV
VLBBNjkfS4eW9esm0jBsNRPWr4au/ihWvdJTlHqJnvPu0oxKEX8J1VIniOMS8vvS
z2ElisdHVsJU0bwcC/tyLBaIMRQZUrDkpsqB+xDEvSOP9FbMbB8lUSfi4BNA1Mc6
wIjrSz/aHH9dZrPMyT892yO+3yaz2WXiPIBF/MrmPc9ere9sNg2Aqw160Xjrw6cZ
i9i6LJnSbi4c4SdHo8uRG70yojqiV9/oZH+oJRFzOjE3+idzpENUsTrh3QorenRw
QvgiONYcmlMS+Bg8tfvH0Mx3z6FEZIIa+kjliV01cY4Xt6PE1bpbDEjCHxYDdZoF
U/O/9bqy0SzPAm6ftr8RxaHEpun9nQPMZqe+RZKfiZWivEZln1HqWhoC3UwnFzNG
qktfNkYmrwzY94SwzOld+yqtnHBURB57dWf+nlpfXiOiUH/FhtzL22q3GLZwfFMP
50v73CnG7n2JSyHhlvXjoSj6v2xe/FKaFll0Af9JkyXn3F975CCVrP587UHVztLS
1nWReSFdW8qwTpuk1skyIMSg2ddQUYsZdRc08jHw1hqkTu8BmEimNbwRo2skw2Wl
QpG7LdugRkca9VGHtMGMv693gvY1quEs2kBEVCQkNue5H2KoGk/MXbIfYEgHXbfu
7OIBKRk33zfJ0ptBBGyCVnyFIp8M5gnLK4azNmluai2EK8sLlWlM0G5EmExKmGmh
/ZVJ4pWPHQohY7hOE0Mn2qpSd77nLTEVmTcLpi7BEo+O362GKuS7co3ZBEbISu+y
c7PofUpYXuLOLcgTcYwnYIAWpsQ5PYPtEA29i5B6XfIeRGHZU2nE+wKoNrXz3Ne4
1UoC6Sbz8nOjvPrK7N6XQkjason0X9+KmLSguobLSBQtDtmocWPlP+r4VKhXI3Pk
iMou0ZlkZoizT3Mh1JxZA6DLU+O20/UYFeYkLGcXpxGkqvVO8JdHWFgXyURzLif/
WhFfPbgjFKEJUt4IOrPsdAUMieJgtsUK2WgE+mMS/WEMooXXQveKAAeWfWossp+m
OKUlTfTz8zWYR0aLFugDndd1c8a7gx6Va/R134+wH7+g8Aj7Rl+GIKDVv6aFuaPz
BgnPVbIUTNyfNLbcAInlKjwhsEF7Ys/crnodTcd0g8UC8evj/smgiKihUO2U2d2y
WK542f4USY9LXCVQ4m+buLBXPJw0uA+6ZWPSpy/KB3nItoEGERm20Hatnb6EYUbl
yPUbQBFvTcIor9jtDOtkQBgo/53YAM0Ev3MoMI7SGgEnpL0bkIOmRgT7H/k9kwR/
Wecwev/V2BgTxjbfZ7Z5dSzUpd85KlNFzbDAbqqPPN1yOnwv28RBwkEgIuNm7O0S
I7StBFbpd/ELTMczRohCJ72YK7kde9+aM+kEW14MmX/4UTsbn0SbboxHtINuRBn7
07TKjpWr9ULqD5WjyOQ0rwE/AofEnQHRsuB/+tN2dwtWtc72/Z+HsKfWlPpacDJl
61HqaWib6WNra/WC+e0PS/KRX57KO4Ibnma5wl8CF4CWc3OH2+0rZ/60GfbVNePX
DnXM1OdXuQYbq31W7YQA6HhEPb80oeO6g1IwjYW2tQ74HL4lmVtqDfJ/7SMpS+Ja
PpO7tzs++ETu9DxlM9vuQYAFwE7NhDwmGNyFCDtoW0dThgM1tlzq+L9ZepWjuWyk
FEToV21GmPV1ENN/kJDl5XPMPM3zj7CZ0sgO4ijRVLGGUNG1oeHFcblxncstANPP
fXkF3APquSBX7O8cuwCSejdT1Uolz3IM5CTN9cylxiDdz7JCv6i0ghSme6++KaTj
5KsqcVAUC7kffstq8/8BzWaXwOKDSA1k/+RjencrpVwEF9wI0/gjoOWKYAz0xNMZ
sqpKPeLhHPrEjEImocLqe7wqFSxrmrvKlhIttyV8F9XF/fa0Ec8yOapmgbh01u94
5rs4CVtEfZSVtcBD9+D1goPeMF208OtAIWC+Hh3ADZwoYf80cAxzVddZ9Mpzv/0x
v7CwR7uW4Tfmfzmnx2MYKhtPGp06m3+Q65aEcsDshoFA4Za1216IdyePPYSQAX3f
X+1SRSm5ENZs9zQ7TnoGRCwhPltuGxvQmoB1AHiW8cmrIldDP6FleEr2Whwv5GT0
XbZmv7KgjpTkC6M3TrGdzMqWKC1XcW6oNHw5gGdw0st8hiBaJZzwPYH+xgO8Yz8N
c99ar/NSwM2r+D188w0UhuWGqNawlJ5f5o+2YGIQqgPP1Vq9gQG0ai3lpM2rfqTh
RSNT6o+bmbhr2HONcRjGkP0dEEwJTcWM0Iotnw86rqs3m21rTmfnTNfpv8tnbAz5
gfWSGLpjC4rBpiQzkQXstVJoN55bqMy3OrGAwpSPd80Ag28wZBCzdzpYt9i2C/3A
J8yaFSXIQgKLCWLoy386G0Pq1Z7afGAUZfwwndY/m4VhYKMzcpwUo7ueguZfu7j/
IMAdvlHIMs4VQsM4AppMZUtucjx7656fPhSAhkhrJxTKk5ty9wdDZK9C7fXWxLMM
/MkK+obD+VBbmqSkDQ1OhMh5NnBSlzZ+vWuO0UvOHu87FCMKORH2xkMkpoJCKpiB
6ZForA3m8G7CQQxsACKst5Gw1csOd9lPcgRpXoKNn1ugWvUgrErkPCZlB6kM2u7R
bX33CfhYdYvunuTOX3ybyrhkhOvOcaYbvwT1LHziQ0yY+bd6ZsXTEW9nEQuTTiNP
RNf+Zl8m0nUT1RDpeJTRpJaNIH14tUjkQlq9Kbeo+bQDqpHcgHWWPI1vk+MJx1W4
WjxEEOod/2vZXAs9SA6ySQCMwG56srJurRMwc78+8iralfUJ5os1RZNrQdBmSWXR
thVRlsyWevrQHEvDPG44Wnv64dUA9K+uJ8P+QhxmQC5kPootcBKeaCY0cSMPaD1C
tOCooD3jCpQib8GgXn2DVD/iKrd7JPQkdhdqA+BYdQE8E1D2qmweuJUh//g+Grns
0N75bMxFPx39WNK0QEvUwkGvR7my+O+vX8SNnGW7L2CkXbpsQHApE19a8NRbTJlu
ZUsF2yAnew1vxe+XdCnQan6gzBc2gMZMWR/ozttL2NyQrPHnciE+5oPzguLaFlUg
3xWCwTlpynPIvHXnMBPOb4Snlkl4FuIybKcYRoCYfRP2p4zfck4fI0RusmdbNR8w
m8YI/c3b5Oz4xYIiaAaTofAren78pw6q+j49KxW2968WXB7G4fvgRvIQQ7ccE4FR
EFMJ1M7hmO4ApK1DOxd60HWqcPNFqNBzjutnb9GLE/eTr0JC5MiCJIdMVxCF3Z3t
UZXHmnU5VYhDGenOtJ1d16J+wTKX72vPtMi4cRPoP0mLr9E3QdSaQZa/8ry5C+av
mpjfy0RBqT38bMHPyFs75/9XznDXBLG4z2QK8kuAeYf4nvpjUCz+sjYah3I/Tydf
NhNTtGyPBQlICxF1kdfq0zojmrm3QwLlW2NNHl+oDjSGa3qjlhS2YdK8HtRHzxPY
TCRpzJeTdl3fb2zR4JTzOWmpDmtmaFLMzbSqPMN6GMdYYquanyS8ERJ7bbGMlyQO
WaRgIYB9y7OGW54UAQmgLMK/6DNXhvmoVWWQpL0Czdk1m6mKNvpLfznUqWZfHfhZ
1yzocthEyb9cE7+GS1C1w6He5Y8V2TtExoGZIXwDcXEHxsL+a7HsYjQWx/w+oIkL
KYbsYuBXXJ7pTLU4ZdrU4LjGnRm1eaMxvlNg+VsCxucSKOnrEJwVYqf/pb8Yk0hs
w9DFzcH67WF216sLHPPn6foND8uM7RuX6g2YDTvfHcu+tLhY444TeKfvh5aQpMCB
rFhUARXoqNTWA5fjSRn/upIF31tBz5Pwwsflz6f20qty0ruuFsUpDEa5bv/K2p+f
ZRpr6IZc/rwC/E2U01Tsp/Mqc5kiWQ7R9KesbMKTX+mgMLxSaeaUTTjoH31Kqkyw
HVKSdP6o48VcYcaTCUZIWBqgG+qv0igPHm25VkOej/2unjxwkfhgAGJhSCMACqe/
rEV4fo9jibTX25VA5/28rw7vFSI6NeH0X0dKXYjfsusw9sglSJpdsDars1B3qQ0U
fMsZ6bEmzvf+Ze1proxHPaAdtYcluan0LOhAxEv8k9vp7tD7IJBv7bTU2WdwzchG
Zz9ASgA6XZfScMS1e+skZBqRjQRPJ5kKT3xOLdVUWoOfJbGOwzJasIdAzrhavBri
gvcdaXji5CeHYrQD/aEeNHN2JbM77cnkfhh65y+okjLKqAUEUYca7vQ1adA1iZ9z
rmEPm1QTKu1oZ9SvnLUuqcvuIxG3gYHskMz2xz6QcDSLdxs4TZ8kPLql39uhtfg7
ma2IXmRnFF76NXzdgfHWoiT0lgTKudurZzHiSQL+g/YGzm1LMUSXKeBz8ukjs2KK
EAhjD4KcVDCTZq9xOX00YouP+WBT5IsrB1f/nUe2KPIucxq6taPdnDQMCBbBWfzi
GobEcOILWeHiGdb0o/NIlv+hl2FAZH23KCT2GzgjtLeFn23IfprOI4OL4Jgx8PGU
RO7tr2biD5J06dUowr+4q/CIOcB7mBgGiC+DRbTIU4jcadV9dDq6cJqvHG0ACWT7
lp7WjqsnhCtULbwUmr4VPaovyCmutRlJdVmGJ+hxO7qUfCdU90+cFBlLlmLGI1nC
nIYPOzQfTTMlVd4e2a+H2Zq4DVMRKlekNRpE3QWccnw7W2jbP5rRDcY0XXoW7xSR
mU21CXh4XqT534EmA20ldQD62B+4Qv5BKmkw0KfWrdGGPg13SdcNbqQOygZOrcP7
Ug8iFWyQOo8NFBNwtj9461fG7FLhaOwPNqB41b8LiBVhZxtFvXUx5x9y5GTJ8tw3
RJu/SuymGMllCeYUW7zvUkug6y13UfYliR+SdNpxo5oAtz6zm/bY98tS/QvNqxvU
1iALQ5X9gvNkVOkuY4aLIhpRxWKgp4kAW00Kk7efmCKNefNaW4GebUYVwD1xgosp
zE2fBdRUf2bO61FrdF6GKDObr6ziznQFkRIHzTs5GjqMZxndeWdCVSWRM1yJqfSX
4W6owo49xcYtGMB1hNu8XQ9Gcsu675h3R+XbtpSmCtTjmXTRHH7hV6G3ovPf2kSK
yrchYgPTQuXKkGovEg/XFWJtMrzqGBcpuc1Y0ayA1WYFj9j8to1q1dwkgSxZXp2e
HeRK0OAuHeorKV4R9cFG5rXp/wpHfSCxVDavEJ/2iXLAwQM6Gu3MYViewkUDcUL1
a3cgnrSqbuPOs07e4yjlXch2fMuooKtf6cvosgpFDfBqgdjR0YCJbBAQQJmTBwTQ
6Ge8KSQbco1FE1JlPLYhf48kXaI7sp6gsko0iS2R1bFN98bOvvp5pK5Y0R4abBuD
x/3+aqtLG9i02GRTDo1kgk/yKN7jjHFnR5CJALx1UL4Keny4H3bOTTlDldaZI3mJ
Htfe1nSR8os1owMAoJ05j9BD9Puk3MEt32XNpRpexWSf79PeLU1sbwZvQgfOFpP2
cwC2v2bcIej5vi9sgoA/A+AQMPG90qgOs1OR9tW2FedpKoM7JTvHP5vWScyz05pH
Nb7F2N7fg2Bw4c5sXoJ7pjzEq2Xx8EgEnin4BvzM1PLHR47pUqsj0k1b7DS65Jnn
bA/KtnP5hOPINHLhdlveG0kxJ9mROF354tONJxkBolF1OpDVXmveBCB2NsIJHM6F
ewkshI7OY8aYyC/oEvjUTjCEbZ0fOsPqiK0M/nFTR90aPpnBHHSAg+XV4LWi8rfc
qM/YpAEyKhUy2oc9tuBsSP43vYhEb5svm4tEXo7SKgQMLsBpbNKloKS2UCWHU/B1
oxbjB70cCCN8kWZ5Wg21nMzZvXHYvO5QshYyzSGY5f3Q/6a7T3rz4zaoilNHEdSR
MEYVbQvFCbOuM5li4y4V/PX9woLmtrNb494gjGqBOXBkVL8ezIdqAhyAEeT1bzl9
AWPL5wT2aUri9GVro+4ETbZGoPQ/Lh98eeduePw8k7u97ytg3jR2zgn+IZ1v2zau
1w5nxML1qcgR4b5ltUcg8eGp9xuGygWR+x+sDfj4rPRgIjRoriADTyiGHJ6gPgb1
2PzA2lkJNz63dUrSy+YUZO8Aq2+IkkBHRAP7BgMwNNH+2cKckdLeLxh4g1+0ctYa
W9qaAWGfuRkzjz49V9NVBJ1CslCL2wXGfk/ioLpRmTieXj56wzD8IICGpGMU1DeX
TRT2+gzpPnx1A907UZlMBoei1VJ0NCocvKnPZ/9OtZ6D3d1hKy8/2HRbzHaUf4v8
puGXTby+a45csgsn9m9a71nzupvp5UCJ37JW2KtKgILQ6fg/yIzpD3S05DlNm+yz
TYUGB+ITc0fTU/4/Zu7paEW/cti3vvP65btwxSDgmh3sY+qwzg6T+ntlNlB5BQbz
U2pzOIvqBsG/5Vt3OmQxIV/NwhMi5Oo1MuxPYUCr9tZ48W2HlUS27stoopHKnJGY
9jH0cywQqjvPrVeN9GoxA1mocNG7Kbq/E1sqUeCsYKi2tqGHTRI9PGYgB22Ab/tZ
Za3EiWN9GUQ6eldT0pAWCV+0NshqH2/cMJXhvSVRweJx133qgiVxyQdiVuM7U+MB
IAbLc6eUSvtMnC72RBPkEGaEYcJuVUI34RJJ0UcerMzu2UpfTb5opHbtUyR86+/v
PMJmCEvWm6qKsoReyyyidGx1q7zpm7oy+L1JlsB+RK19MKVtvCOVV1IwYN8KM1Sg
T3GP90WgQjXCOxbqdJRPWxswXAXehQM+CnAUN6SWp2rQILqjpzAAQrtcYFyA56EZ
qulJ9QGE48bxq9+7MG8RPxc83Wvcpbm/gfYD0eBfntXQzw0cD+2BbKZBjNL08B7/
EPQ4hjXZz7LYgFysAbEdj4bj/p7wjw7dv6GRQabMAqytHW13oFYjywD06fhugifR
Xl4IQ9gzyikCFMICKmod94jCtbxq19TKLSzoEGU3UVFbcQO8UgS81MmPHOR8KMjj
4vRphupB6Bm5woc7yHk7nnsVO9XFb9TGfuco7E0PIWkAMpPOX1QwmelP1eA0UZnK
agPdi6BcZJBKnQN+bNEBF7ETz2rpxcDmp6IixH/Gx3nglUuwv65mxo8U5wsNARHA
4cYK5MDy1WXsYToYQ9d24PD8ePwvddnwl4hCj7ijpcxghmJ8zvAn9HcVr/m520HL
DhtxxaUHAHa1SJkzG/TkcNxMNRqTCsoX1xWeENbHfI90hCD+9tQEyaO1Q6Rg9RwH
0Aq98YWPv6XZSg2Wdz7D8G5M4oPuUJz2jNAr6BdZ5vyXAIISbCnQHK0WVDqCXTgG
RgmSu0Q3UUXsqZM+WkdJ7wFFWkB1Vn/jS6zxsuW/RVUJdOiNmJKQYjuuJifjJWAG
EZChNn5oesVvssEyQV+kOzRUtgUEYiZiP3YP56mdx5IuXB9rrCQOS0dR7okZYd1+
iZ3L7+0fAg62DxE+OAS4nR4+Mmqw7UDVq6jLH5EE5tWVg9FIwLHyLZA9L14zSSoM
6DKa/bushqZBymqbqQPtzEEXpkXoGbRiRld/FYpz2Ja/nb0i33xW8Y8KJEdMZBPu
QnerdyfIw3uQoo4MKbo1EC14/FzZkxl4ZVxgahvLeJ1YysQQGhA2mo35nLDfJ+tt
ffIMz/ZVbmy627beDlGHYtnob2cEU7go0Ag6jea6b2dHhyq2i8vrxsRPXziRpEl+
X5iya2he7PC+0rrVNmeYrNEWhQiYgLe6silycVxPhRbgyLn84UfsVB72Rna+eXI3
aHpt6A1QXNELveG5vt1ZixbsoO/QdAMfObJyumx+JVCdzr/YlSRIYZI+BItvI5TM
8hCU7lsmf463v+DBwv7ew5F1SuJn+2cg+dhqaVSCzsgG6BO2tdBMXmnmTvSCrsVO
xzDuhAEGZxa+VhhNkSq6N0CVPnfJezc0ju+fKVaVeFNjOYTC8NW6C7rAImjPaG31
CVTiUnxXA/ReTKB8AaB2i6GWbe8ppDlzKjHOQuDHMW33uu7ELPBfTiXD6MZHSt8d
RraobmEA5Z8SbSvDRUCVBxd1djuqqj8/qLgYw3JBYCYQ/j8ltm9OSrIukWbV0uXA
aMh6PamaQtxRsquHvWoUpIoTHOzhsts9tB1mtvWdEm+mIQlq3uYIRE7FVK9l5IQE
nJBqqAv0kdFNRB7adRgy0pMIiar8COGp6o4BYTSN1hzLcqbcb3BSPbmi0EAfza0B
mqGGkiHDp8llwOgpD276jSZwhEEJ6U7a73pdD5mHBper2dTSuGwtN5vhjLBtZ0b/
UqpL2YT26Xdu4D7G2ErQbZLThn0gKNZmgMRjgPptSzyLeqasoPNkBTSVbU2Zq2my
wWk8DzG1CqkfvjO5BV6eDZCL6ymDBUR5TIbBKuxHyr+zFfK3ojPYckYJnF1z1Eyv
Y9bzvrowscYSxz/7sVDu+O/Y/uFQ1RBko5n4QcyyX1sym2KBuBRw2X8+fAKuP1qe
fFJLeMpeNd3X/xK7IYN0ffZio1+ClFCZ43j2D6aRvlqDJ0i08rXni5sx2WqWrRFj
agNYZts5YI5/cg39+W09T9f7Zff1eBJ9Of8LFclHgqY5VhGpn4oInohWvxtOJvjM
SAQRM0FoI8MKMDjsLkLKyX/IuEecDknIPQ5y8exyMFT5YsZAe9Sw8gHRShU3y9kX
xsZtXhu4ujNMTKw0073VPxaYuwAmZaUSnpT+Dwo1H9abXHqMakR+w04sayPESi9X
qjzAKprTikmgUDFVGH+qjCvM1loPteVpkmNq5VCO1mX4cRQlJZx4r5tlp4T8Q5Bq
vATQ/kaULw2lO08IuzpwO8hFfAeiB9NFYNr+oHCIQFU6q6EDXFzpeFJZanPKZvzf
uHliAHxpPvesUwM5ev03I4NrXH/zPQ7F8NyKFa45/pbT7w7BqN7UEftNn0IW9U6Z
oMy0HsVsN9Wk9SToK7Mt1VhTQeYfsVjBsH57lVeRdfUM1AExKdymyFPRWy9EW6/v
+KnwpOhFu6tmGaz40ZmMgfrc6fRx0n6CfqkgZKuwk1G0d74PxspSrCbY+jl0QAni
ZlrJUcM4fquFgC2m+rJbDW3+Pa7E1ggm1YjxJlrdPSmQ0T1LsSwZHcsn94neFr8q
Cy4MFYbv0VCHfrUT7eO2ah82+GK3H5h8uQLJGKfwshhOjFuUBnlkZO6MOAc0hFWi
iULGDaZ84CH1M1XfJlS357rZYaLRcTUzwGrj/iHO3faLSxJC0ksg4aAUIESjriqW
KIqWA0X5tKcchd4fiqlELODYIRxKFHOB/bstsp+3GPgGOYN+RYwMvVULI9hJqGzP
hfevpKZm3UY6K1wrY5iEJodtm0Hk7nRybzluKtYr8QQXebG8vI46bhTGNHfmySg8
3NGQsZ/7lEo7F/H5+IL8ladiUNICcaLOiBN+lhUxu6ZHx4pf9skF91mrTv3WZ3Oy
v50V7PNPELj5ua2duxw3zEQR5eFEBjXt2KbcedBh9+g8/26o3OZxSfuxdrFeKGT8
S33YJ+LR6szvVFJ6SyWybQ1rRJ7MFqpJPgtudMBGbBzBpbySK/oKQ6k+3MzR8Fm0
X2QJHmZ5IZdCFNnbnc0x/eWFADN4o494mw7YLlowNHeEpmOZH/PmqbARfc/NvHop
gbOWKvzsYccISDqssvRWZdws9QgP5LOu9sBrlIeOzIIKycKwxCA9ba4TMOdl7aJL
Qj9YfqMy53fqvrsXSN0jxM12lTSMgUBP6oG/OnZorqkc68DxTkEFyIFJLGJxhMgi
F/nfriDRnwzeDGB66J6XT6MngSSEG6SOBLq/cEd1u7mjeJRvQgfTIVN5KI1RtSTL
s+077krme6GgF3jmu5HO26THwq1n9pIJ1paDJULp3kbEqcwVKc6M+CiUpmao4vpY
htz3oIiemSuqYS8hYWE8hYEkzhUQeU1u3mnoEA8dyHxurhjYPEEDw/jVnLSOx4td
mlNj5Fcl7yGu0gNTtzKrque6mbdT56nDKaVB26F69QSYb4rwPTAq3JXoNj8zfUE5
Zu8YvRNlc4Mjp9DeAOssrlJ2nFb1/qyi8i8dfnoW7NnpnQt5cG9wXu0392KpkbIT
OjbEGFIJ3jBwG38m9XkSgbD8eNJzxGO0ulaOQxgV1AlPd3zjn27i/8m+O2rJwAjf
yqJl/zXLQaHBUZd82vORt/3ZNom8km6461SeNmyNNYBW9WEYYRnKLPscDTm9hK2Z
MbDNXFLph9pO1Vy1o6L3FvrfUe/t4WbfSEvFYwbj1na3T8/aNzzYUMy+qNjmcQ+T
wWZcU9aQYA7RTiT5qLZvBwsNYvI2kkV2CRwRfcrOI6lqgCDdPNKeKsyBkFOddhUw
rpF4i+eFB5jglYbND6poKVwk7PcmwOjlO0Zhgjdp2KixeBFcpUm+gTcOUYjPISs2
z4O52yAdR9blmEpkXWv/8w6/3W2vc4B2149/0FOpR8IwqHej+53xYk/fDMZ+fW3G
pfno67bIDR9f4vpjwr0ArS12l5W5sxXPiCIW+w3jWpXCy17LubCg/PE8GymdxnkF
FUdWAik44bRYR1AqIjTVAKY7llpTS1OPJIxiYNqV+PDnuk7qgtFBYDoGA6ZG3AGA
aPE0uEi20O0NQnv4IFRpm8lcwKbXyxnnyUvynBUvXxImLKn2lQWaULxF/fv7OzJJ
Tf+hMHUfNckSW53+H4Oj3bRVeT+rCSEiOfW3+TR7xadi5ZZPnub2Qrqg+T5SfNeU
5oVGdDe3HU9BAHuCcuPI4K4FHGxBhAwibu+KA7wdY7OG9Od0k40Hlavrk/ivM0v0
iEPZKyz0A/Rli7OTPVohsXgTXsuUxEhlSup+5xaFgq9X10fVnktS9oMOmxSQoq7P
uET8DJ5/D2weI59HVX4w6YaQHrgq4CNuIqljefKfHgALfG5aVq0DQDHH53mI4WRG
uatjLyQjj7DRMSSSmw7yGWMadmfLa4CRyTy9xPFH+1lgjn/teLaxvDhj5qaSx183
+4z185/cBNc6/sHnpOLdpqQ3P4xtPhb9tECcr6bAajTtKDvcEoHsjYbGkULtoch7
4XLCMjMO5Z1hFWQdj3VdCLCz2XWYR7Nrjvq52IF67D2ZdPdAJ+g29ANNQMVn6f1G
WJYoyOxEQurMpp/MkxuqgheaeQ4xBEQIVxOpTlEj7XR5Qa22tDfWxW0q+i0P6ZIR
FUYqGjNx8901dgMlvhdJ2c1XigRRXA+s3WTC5O5bJcPfz8Ctawg+8lBnxz7h67H1
cjdroLe5gRULhsNUuFDGi6y5O3t44fPw0qaLmdpu2yRBkiKMjQ9Ww72I1AJb8+Ai
yoAjqRXf0GXmJwkC8n2CUBTu1HjDQRu124IVGcT6JNLHPzCrBrK6+75BGnVOHq77
mmodb1NZDGWYq0SYBSr2dPq7sRQhHJ3ALX8yPVhH6ADmGHybOdTcmwdkiaZZJyrd
XxPg/ALQbkQdyPIj1Bi+XdJ115f77a9Mx0tWr2BBREFgDLvFmcBlNhiVbFsA+Mx1
UrGPll1oe5aBGlp0PPLmtFxh6GfceH9zshxmltQJfk20EU1i6k0ZmtgseYJjA8D6
7fdvHdWNmHDLkpVdPKCo+gwiUhjpgrIniusly1nrvqsdi71yKBKw/yl6q8RlAkjk
z64Unkgbh4tn6lv0t0CvtG6Pxyc8hqScgKsLCBYuc7a4IWJTYNDAtJbA6+haYrpc
AAjIF7C8qn5ZSbFCP74uznaP7YXYGq5ZuGhYdwIjuUZRLWWuqCOIhjy7H9Ey813I
EXB1bt+3h4z7aCMq7UoKsB7xdElgdlSX1nmyuwlDVjy00rVk3RJyK+ERi9fS7VAn
EyjXUTK9jlpQZVq8SIB2p2YGXUjUTJpZUrt1Ql68kkmFnRJIhO6iga5TWv+9Fa0r
I54+rFccvcwnE+nr3g6uAiniaLijfJzP8M9OFWlDMjBZFkbthxG7zPA+zSPoCPnT
lZ+kdGxDuz0xfkOJTRsWkdtha2bQLBSSiq70PBD/p7cjMc7pKh3VNB2IXFVHTeG2
Kyl7fVQA6BBcXwoYiaoKX4dGJa3shkPfO9nq+mzGfhMk8iotxJWWa2LFB/6/xTTR
9skkto/5jqC2LpB+x4POguC2I5MvwpD04yU/UxP3oUHjCNuEZTEe0r0G8++LUWe2
W1ocJ+pzfhWeOoqjkZLhAUa72rZcG2vEHAKlXr06xKF9VZSTb/i+EudHs/hdVI43
BGc+dhYTOJ2/SLoFqvQgp8ymWDsO8DfLhGlnp88MIoDatOSz06WBHYebrPFqv79D
bf2MKC+0HcNQs+6hHc513LcQWwID69kgDGvTt2pJ3ZKQeriBVRfu5iXRG9ahJ87r
RPngWT6dDDtX4qeNwupNN/yOf0HZbnlXEaT5gN2T383GwBVsyxV9g+r+gn5VYvA4
DbHK6NHW9kE1cJnMJpLluSRj7ktrbnh2PRWjBA/X/pILguGKU4T2F8+MfcLAUQk6
nFYT/b8kqQ0DeVxgGqhjeaBBco7coeAwDgVnWFKApfcaLd1SETNN26AGrPrM5OvC
c8Bp8c28Lo7CjfUngtkCd5siwIBxDmpGDnWZKbpi4kl71rR4UeFK+MXHglYTU9Ai
vsnz2LQlzS7f4qRjtKRUdecVo7lAsk73pLRKkp/B5E+w3/gaKJE93J8iA4tE8xBW
SHlXom2CErDCg+B8XIY1yUt4CuB9jaEf2+yJ85oDqXCONev1PmVG4YFLApg9Nm+o
CAaBmZ4YtH5HUbQLcEYyD8VDo3zB6N1Aj2E5viT+CUFZf0z1e6drxFkGbGky9Hmh
nFEn12dxAc5myQ3V1i8w5ApUlacFImOZpSQZ+wscDLtP6kLI6q3FiO/he2UujPPv
i6MyaTxq2GGYb2gN7hImulZYSdlUALkCgf7zDd1XFGeesUkIxTb2etAMWiGM510i
txYedJ00tbY8dar38+yse8OqPWR++aGLaOTkIY6hhIz6z2kaMV11IrcZDx5fcG+N
+aWjH6LBUrxVQmA6/UZmCTbon5+cZrzhTKNKcmaaVgcwsWC5/+3sRBpcuKCgK8/A
4h3rwnH+PHQelZqSCTNSAxWeG+ZkeDQf1QJqusGQbfLYom+lJGpZr2yGJA1wUOV4
/JNr4fcjB5+whFoW/QeC3gIcqTgbzF1mBLsR+3fQtZTlY/QlABaz04yjg87zMJU5
L8FlGLM/TYjik0wRTOBibyRfCnPyu0bjyvlOQWCF/CCJrWrHXNv2ng61gsFPxMuc
qI8QyZUn/y/niMMoNaVqCXD5UoqufiAHhJZhryfxj3e7K65lxIgnxr9Q4NvyPFqc
30tXRtAynau18HGwbUDuUwE/wb8bJEsk2tUSfdxAZozB24v0BLd1H5dpBTzQ9BJY
7xEMb3AaILj2oIb5LICahSd+y7TmdGOG85ys3rloWWSX2Yl7wDDhDUVcbeu37XzM
fA+UnGc3EN5suTQCAxhFMTW/Ov5FRjRDedKgx+LKdiRw2bFWhpRMdiwo9hpvSyp3
/PmlNs1HRR4Llq3oMugrPQbaaK6lNs+C1fZbUlQCioUM86ONPe6mz4jGeEsItiMa
KlPgKbp05FfFeQw1s5SSxHQqrwk/8PLplDMXBmSFyk3IqukdIdb9ptumiKV4Pm/9
TqwtMAQ1zDRjJdqGu1GfGsXMwyIkjy7Jv4klxQZXVHZv9/lmLxVEMi0KbhyOh6QF
R6rSPO6AgqRfFNybx2sPbj3vpJ1dDyQMNm+IB4QaqspKbYJWLmSSJ7cLDadvlbqm
YtBTwtlfCMMktwlA3loTusLYb3bPZCLdcZuptNWKb/jvpGHZaTurNeyFjLS4AqkD
7+KG+ylAF6kFgQVR+Plo+wUX377K8bBrauUwr1Sc0KeLhPkgipHILC6OARl49ZqW
/AvfxIdC9mON3kcNEuTfqtYmPVOL7wstcx92NiYm7WjgMaxTm57RRsmGST5JKWKA
b2SpjaxNpSpP57CD2FqZniSTFh8+DU8mD916PFHJlfFZxI57fedaG8/ZeXc5x4H4
3h61a8Jvq2Ao2XFlDmkwluB4AEipBiGyT0ji+a717XNp253nclfr1AXcmv/72CeN
brH0AtwA9G0+zRHmyuKdM3T+3IAB4xVr3E0JP9xERIMdH+kQMjValfIA7R/KlluO
I03Dx3w2A16T5BdOoVFzDHEyvfjkTfb7W5hBjiS62Bf+gKSRx5sp0MnnbO6m2hhZ
v53/FQNM6QlJlcYh4/V9icbBYpkPP+ePpm3ng54GuwT5e7aglmo1jWV0GFs3KAr0
mo7jPp2gYY5gYa3Bo9s6gd7XnBo2miUiZ8OcV+/kUuHn0wEw0XoK+gmOKAZMRz0o
pN8ljGu/L48EOdHgPhKjz2F/0FBK01/3qkYvlF0n/La8cj5sDjkSt4sn+qYbJRZ5
NX7gTvbABWLPxAiosIg9AUGJKg/SFnPcg2js7/1A1R8egjAjNceM7YP77wmS916F
/6Q5vQ0V8Y2emJp5pq1STAlSxLPKttiPYpy/btdPXPDyxwJtZZZdqyOylr8vgGf0
7T+jKAZLzPZ+vFk6DIlXxUkxjrxhiSB21uwILB9MhjMXQJTI/BrpSEVIZF6WqIpI
fqlxx9HIyStltSoMWZTONqynya8ueX5iryf3+oJrx8+W/N0/loEMh8LSIydXLX1B
HewhKuKwhbEw+tONeB31/P6a2+NmVSCucrSdrWx8XtGTmYM/zGyMrHoaq3Pdokk4
rSciXkWWOeveL6Vabo2rVmz0FEVTrb6/zCcfMw01pUsCpPBvmbv0YnwGudlWFPJ7
13bpvls2AT6AlqrX5J8/d4APFjzZkEqflFlBk+AXT3cPcC52KUEWBjerWG8hOSc+
nLOPMMHq+9leShfM7qIMx6b2Lqb+9p/htwQLxdyPmH/g6kT4iIWWnnFKRDG9FubF
2eiPlgQflRvj04VSi5+reOfGwyTP4JepYv6P4+xEJ+xsl/7Sy51BNHe9LlaPOCr7
56MAJpB1QXGm4ZylFCCld0daAJblHgmt7dKt5sl5xM6Kff8pF3oPXiBWQOY23epn
jNOMJyjddOwLEGXTR2mvrRpByaAg1S4CCf7O4La9bgb601JXS0BWRmRz0fWWCw0l
AYZ9HzTG+mlUVCKLpV/ptm2kmeKZicX93BgiEKFVdU0DunA7RufFlUaPy2KGuLBV
Y3ZIhe64K3G8tRHFjydZUdU35qZ/sfeldb/poo0Oh1l7O6JLsY07WyoSen9j+Om+
OoPDhQEsFttb9mdkXH3m/MKrx8re8KOLjPINUpg4WTRF26UQGKI7NQF50HGvSp2I
XxGdroKcgY/x/OLWYZMw8B/biTcpdN2GTP6+v6WujSpnzw1kwUA98bGMIZqI8sxc
w3pCs4jjHGHEpepVErLRsFvLJ5cCo9XgFQ1GAFlA/oz8LRUYi3lsMN6+lekVrhxy
C/2JZCcw5zCXxqyf5ejyia5Oa0avSQlCEWzUXktLWdrtFNzTmX95RPe4MSR1HTGZ
/LO0FZEnd/mXOO+ItY0zDxRsriv2fEFnbdowA0PXIq+SpWQPzjegZTKW5vTx6K+L
hDMNjvi20uC2sxleAcFgNsS9AH0WFvDU43HGb3iVxkc1Rb92CEeFKRsWP+0zQRbx
fUxsYskEn7jPhOcdllLck5L1s56uNmsOAhtp11LZNPICJjybVwJkeR8j0csv7M4f
V/0/OX0Sh1uy3VETBE4WYn51YhClG4M0ydSU0+6oCQISMaveZcmZYiM/ZNBODvpt
+k1jHBDzduv+qZ1fVdH6Q3hgOGyUl15qCu4Q7AowBYTXgdKEqiLdZLHGte+5eLgD
PlVGeQJtsJqPbVCEbDQfYY2cgtHAzw1lWFxoxrRa/bOQ9dCJZtvqslrAnhApd4z/
ij3rGhSKjyQ3Jjzgcxp9TyTfdBx+M5WYAbW5YYxibTpv1R2sYRsXI1KvXKt+KJAA
cQFE0UYf62LlG1X3lnYQWHNdHtNDsVE+RaYOzF5578hOsUnb4n+pIjlqO+ZmxhPI
laVYcwqlOZO+GWhQwbK8pLaRUR4HbJBhs9jUChqmBbIwobRWQCUrJNAaFZ24aKbv
ZtA3KoNdTPeI1sKkS1Kgmwtk4GgTzZfFSJs2pqxjLcdVAv+CUvbtjfqr3z4XlzUU
4jG4Ua4J76T8SQvlzb6NPgm8k+WeHIFxQX1cMrmZjhPK8/CEzTvzHUf6ImTncscw
FJyW1z4JVRLFDUzJRTViTV3/QiPUaIgX8sHhm0bFcnSG/K09RA3Q0wsxti5RB+RE
LDapYn8iDO9WTLZWpZKu1qo9OlzedesPUnMYPIIXZLI9STh6BS8l/0GTgbZsUbXB
3+xLcT0HPmAVzEuGWzNWfkgNl1RsZ9h/7P29bAo+CZRj88+tVBeaX29Tj3048Ca+
pwy7kJgDTzRk/kOyCmLjGntEWmjHNtT+kS1bSXQnl3KVRXDeLAB0HgS0PvPHvwEL
kV2TMQ4ifBl/f+CnU1wsBwHXsUMniHXJnFjNfudmfadMcK5FNv8E3/IY/8Hr12HE
D6dyM0GDfKjnTRyQJ3P4ZQusrYczDif6s83XrGLq78+OMmL5DqFrW0wdNQ3nhcX7
EZR0ltyK4EQF4xC8SoIdBA/KnbrAtd0zGmpJuqo+peosGF+BeCnStoOsSLUXy8eu
A4pX21T+0RbsdKv2hQZIs3OGfYxGYY65/dC2tFoVNr1D3bOi8YXzLL/BRo1scwty
EhEkyBPHqMKS83EGbpftD4Fq3BQ+JVERW++t3ha9Nw4tYfzi4PcQbcl7JeV2A3ne
fBobhDJKgWjLK7BhJrE4ImcHqWe4j0umixOIRY7SCj/tWV7urWjYQzdX/15FOAsA
ByWG6mhNo4nA5+O6TXGKZbrptlAnBTe48PkGRw8Mi4hjwG5HlTW2nfk86cDZfFEK
8YpfgIpFWrLFpsC0nqC3k4Dn3RaNgFM538EqroSoGCkKsAEquHd545ctA0Df30y9
TYsEAwmREyFOV7nSvwbpFn8bZwLWNgWAgNV+0+M0hBU2Nk3EZUBjyFJMVO/yDHHi
vh367suIMN+GjNVIiBdaEA3oWDH3IGWZ/6Bh/7eLjOBRw0+KdjhoDlMmCOh2bDaF
ydt+qa87fBLKxsFnrCCo5x9C4RVWL+9QoboP8NTeod5ohztKuuzW3BVURRZU5O30
ycINBXsfP7zibKvIo9H+T4SIEYxpjQ+SRkR3CITtCnKvkXHesKYpYvBqij6u59vR
AdE0rCze/BLKEH5k+PgeFFXiftWPbA0/iFqrkUOx1H4Na8b905zvA1+gSgrnfcmm
h541W/PMOpxq/Sl2nF8RUAzq/Vab9q6XtziyRXKBw3KbzT/G3rDXQNbv9OM6WRDe
76Iu5f412S5yiJ65QUEJKQe2UgwCdSsb40gFEuzCuwc68tSTC2zllvbqI39oHm15
ydTe87V3G0bBR1qM7JdRWsm9cPu/6rujzT+vS77CSgdccEg7Mw1GDjlRFsMUsGHF
zGVt0irnfx3Rj/Qg+ZCGsUZoIR+ceuBugo3wabRIwJKyF/k2rVc13geKfMnwCDmI
HzcBgDd+0Tm0iLXYnQ04O2mM7kVsuCQyys5lEzy1IOGPyuO4NfeLvLli16BsSuk2
3BV9uG0qyaKf2w2nk1cnE0wV3oci0A4oD8IBXpw2kaJlCuS8Na/zYuokzRpxd7pG
Ie1ROpqNSey2SnMKrSUTKonpGyWR8olx01RA/ELNbsiHFekwe7AyIx4dUr9FbAlN
ytk/qE5nA/dy2X+vMnbe7jQnrfLsviGwfY01uOlaJHzrNNLmZQsAURhfe5e/7rVs
0sCyTObqP8FQy2bvpTOU2qJCBgUIaRDNmpXD/80vazxLCnVo7fe4YWXnhBNAI/CB
hr0xus5OpIfiECmZhQuZN/3rbO4rmJrgKkNrLbV8NAWNacPWxfBuyUJJ8l9YneWh
NxG4RiSaVr5Zm8/EOdOgYX+Wf6adbi8DWW7iObQviM9M98SJlLN3Hlmc4lKuuoZK
80vG9gDnACOvAOYJklN1qpJgMGBAomodo4W1XBr4z1JjBu36kPHtqCAmIFglYZll
I8/DLYig4jJxq3bOh7kJVJi0/+qWScH0K8oOoCeW6Dza/NQG9Xspv4v6BP/YmDbv
DL3I5AnduIcRHqxg4gj6sRXGy8Dn90J5MxTxEeVYxfJrMzPHDkyCbxZCLJbzE/+S
77ZUIt50oHxZX+LDnONSsA2rfuEL6Ys6h+cRGC1WkgT0DlIk1Sgp6Vsdmo1yMrL6
jnrJ6FPUXQe9FFe736Kd/2vuz0tC40YrJeJYOQvwzuAEd1FVLu6sSJMnU/7LD8ss
j1zEikCa02TC949ewCU02vd90ZcDoasinJRuUvCK/3UF0kqZa4x/G66fUPIgPQ2b
ua5qUPAHChowqb+olWVgc+zcFB7VUxkV61cYA//QA0l7AOVCBEAJ0w9T2jvtf8Dv
KcXd5+xaV1I49ERv6KgZYb+eeD0MN06OnusIKyA80j4IQKZ+t9cr9SDGQLggrt9s
tYjMyoLfh7K0bgygZfLOEuCY4787a8Nmoog1BOpi9DJ8GmvyZdVSufPn87oIpeB3
Yz1RH2sVmhm/FxHbc52WNKS7970uBF4o0v/DTdpZ2kXaFKpwgyY8ALeXVzihQEJN
criUHxgT5AATlExi9hVUD3+UJBrlgpfOtMQWpIHwUY5UenBpInwV4ScfvViDCucp
kNZVofX/DSBb+jfp2+t89dDcsNroAT/KcrTiVQLHFiUd/sQxWdbYFaHWpDcGmz+A
SN2qTgbs4jxRoMqSQliQA9a1tT2JN6CL8DmifzgKunwglR3XGH/J3yrKlFp6o/v6
l2HRm89Zo6ThJCjjr/SQHsujf7jnPS6LuMVOLD2vE2F6x2aFyJBe638MxogfkXTe
3Kpf+lnbk80opkwqVV1secnYw1kEojUh4gSW/Vsk0YByFZX530bEhwSSPQGp8Mbo
6zT3YtkMVKGTHbQAm6gIJgZNMgx0xg0+af1XAFof02LVrfLNPOS44opj+AhF5Hmi
S04SHRycktw+aUjq1otCMwbo2B0SkIjASHCkjQ333AUPJ5o18LcmttpN7snIoDQ7
1etg0ldzgQxyJZ7frV8rQgnnxhYaWoOdrbsN7/7L6YLfSztts+JiPDtt+vaDcjCq
4eo4kRhGKG2zZuIPtSJ0cHZKIaMoB1PGfP0F7Dn0UrGTtkKZ0P/v/T+gNqQ6jlEt
pDjNRu8BP0n7V715AdMVrpHzGMWUOMJnfFNHK7+fvSHQJJu6XAVyxz0FuGnO/l5y
b1fZkzaIqjaYcupDmTN7hk0YhSg/CsyWRN/Nb1umw41+rrpDicfWMyQ69hOEPH2l
L/z9VugOI4+QLSLF2CXmsUNQjvFgBd0FybDF4yBMloQRWhT5YnDR8GsoSq+X+doY
84voEdotxn3pmx8Z4FdSk9ha7DEhaD4cuX7A5doSSWujP1TLHg3IgPesbyFzIAfJ
IxNWpl4qXmvBnoGomOVpxNM2m1vrU4DnsC6HFhK3vp20EqosKSeiruoGOr+l82KX
ZDN+4FBmE0Q3QhYDMNSTyXywfTu5I8G9XX4c+qbo3taO37QNpE45J4j0g2AxYu69
rwTV+5QcDCBOiARbj17LzkiA0wTVidl7eW3xTsGC7r1UKMQSYl2zob0eKP6EsVmB
rd0BKBaMn7EwXJREQnL0NpiAq0SyGIGCtj7tvcmj5ze6rYtALdAr3NWAEYGE+Y1o
SAhR3V4PzTRd5iPP/pZ0fLU5cYd0hujtAGLccTfFKfctkox2hl9QadNxCoC/emev
plhBb1kbd2+hi3ne/riEOa697C1Mlwwg7VDrWsklAxFGSc5sXwuCdMmULbXRkjLh
5g/JukauEwpwwrynIYzsjlOJd85uPEgSN1xhlZG5z2mfxy/D16vdSAHqBoy9O4kz
ExeN31Y68MBRztrpMYgnYII4ySfldINVAtTDLKSPvO0EII/ojypOQwF+jyTqpwGh
bV9yjoggFWswxyJ6n2dn5zfbB6x/bHRQaZpVVgIjUBRWqZNi1P0NuFVkAJBW4jiH
PsyhnNWXtTYgGSgQSO1gYakLaB/9jJJ/9WuVAF7x5XZdxw+KYxVI/XxjOH3BbjS2
JuVu1lrbaj3e9OID5dYgmuVVdG9EJMGYvZa93loz8O800BxmzFdMX57sIAaP8tfC
cOkxuqC9XE8bbYNEBE9cqJYy0+fdeihgQTm5IcTsWndr0AdEPtjFsIngIM3dGA7T
CzClQGPpzNgtsbmsPAexIKR2wKPch6zv7BKvumSZ44rv+kpzS79jDiZbcQ8zR1Wp
1G2wa4ibks+KoxKjfKh92Vv7QkOH6oslnZZwisGMp1d/8SvMTAa7xUpiJFGRQ35g
iYUMLhwkzxqmoQibLJ3/1le+cxLKcD0AnNuys9ArgGyQrWNQnvNwGpoXI7Ve3kD5
02tMbHSx5s8senQomkq1wGEjkrRgI++iuQYD+XBgEzDwTR7Sz1n7zFMihlXZyT+3
YxUlHY40xbrmR10awUTR6Ch8sWvgFFSKIYiRRSDaPK6Pxmds0JxOVpnnnKSXpKXk
Zf9fel7h3hpZD7mld3SlUhdvQX/J1eXcVjTb7lVuHbnt+p7RDkmjD1fD+yhTO6VJ
ov/dzGNfnHOwiIB84OYwcPcRqNZMIPxnXao9xuH/FPsHtwn7fyjGBDiJdSh794tT
3M2xtZZEd/86gF4U1dEu9AP+PCsNeQwPvdiW41x0k0V3Tm1Tj2v+FzuKdwRKCZNy
6S7kxEZubDioQ6UBxSRQQGO1Q5fcrXjjhGLq9K3v8wKxuk2FyTiUlwC3fbakObUj
MPdBLygP2Sn47Q4HHD7hRo7AkCPkIytiWAuwqmtVgtU8kJzuWCqLaU3s80XNwO13
ZwkvwXCnDk2NYaacV/HMY2KybPKm7C72emCWcdo/7pN5tN8H7kXTBDfNVxjViOjU
pzfqq1YzmYXZelr4Oj1DSZJnAwgaN7wkMm0O4rphVSg5hI1KXv9xPuKN30uPBEna
U+7p4I+REo7sR8PbHnqfExAYaVlKz7QHhieFuYgDAYXnB8njPgRuNBV6TnSp6rwB
ST6tgy0qRZZNn3nLe12hGaW8BqGORePFzlBxCgUtLGbENg+A8EJZ9dTkMGNGeoos
rqEgXl14azfxT8Avzz1vqmlHzA1J3NiPRhwmNUrQnzQOKU5uwDtKq29xqPaYcoV/
ojKQ7yh1IkWVsNF+34QtTKZql/cs6LWss7nVNK7sQu9yE5PLxnp8D/sfIpPyJMiC
Znbp1vqyJw9GmgN8ZnaBYLqZ8DJZCgF0V74duvKwjDuGpUZ/VfI6E07igDIDUm9p
7eOlvlt0SRBxYE4WAl/A9GNrm7VqKP0LvkDZoKoDJfDpmZ7wRLtPGkGJDa64eJLr
keBNmnm+Kax7H/DiPkGH4rEO3JLhQ88BmX78V9qRQGS19xEiPGQbnnkk0A13UopO
Ui8CmpFG7VnYLC6wfvzmoFDqknGX03RmHzSlJAOD7Yb5sn2SptKyB4RArzkjOngT
hkGVFkQ1AxUdAQ5ftjwXKfmo8OYGhMxLKkFdaAw9iIbdohPXd5gO/0H9f1v7pPc8
3Jgb27uKgvwfSzrKhbOIAgxFJy71lY06uGhu+wTfXOAyZNJhxiNTWvFlp9lB4sOT
mqxq75skzhq6lFCsKR+VJ2xE4JI1BlUFGIlim74x9dQDWpYXEYruLqM08SBMqBAU
rmVuFdoALyCVWyUYWkfHmGfNK0ZqaT+vHTuUOqMO/mCj5djP/VCdlr60OtT6sNX4
YXQCsTLyvs6X5eXk28Uwkqvq7b1wGg4+w5EGiEyX9wEoTfwH+PI/EEBPA8MevqeO
sm103OOTF1GLGm18xuHFa3MWzWWwA3HEjhZx5eky2WQN/bU6cFpnmNBuasozRPuq
0rNYOaaJDt4xaoCfWbrCmIDz29sXxR0DWxgzJLnZVz1Yar4qy89MH0StPvIhJvPs
ceX/+5BBITFQ/IFZKmodL9YTVk3fjkyG6jXqlfJh5YEFdgrgw5wngkjeMGOTG9Rp
8dgHR1/8uZKRzginu+1xyeCXnRjchdVwEmu/FdQNFKMkRr7cV9flqU46pg0tx1WY
J4rt7qlO/ExB3eAyd/JDpheo/AQvkcQsqcfxf/lgumk+gS2TJRramHFm+sBfDdhN
QXHkkdLqdzJjZDYCLRm7vlJPIjeSTkjVasj38zvcWL6RwVIgsK0bnkTrrGonHcvi
wAhfbAym4Z7c6PxrloS9QjFnIzN4HWFHchHyohHS3QbO6K4JzUM2RmO2NLVRUim2
awvvSoG8vZvdtnKv4WGaF7OoUQHTKi+3tYJ5enPPPlCLj3Zv1ceCgjT+5GqVLGca
iddI+PJCs93odfN1QOUqjtmx5URkrE8n6VF3s3Q6UeFenN2PCGcICCzRBiPjIlD3
Owm2I4vkc78t6Ss42pDd8UetSx3yyKroR+XBML9VwL+zskBS387xrIYnzfREaoIX
EqS2YpvC2v/smH8YFq35/wMSuVSA8ks1WYE+U8VBCV6MBfyaSozrzD+owmxnw0Ss
VkC7QwP+kY2RvNrxkioQO6AKhG+c+DtTlVV33yXwNufVsQqSkJ2saG5eHsPB/H30
k18kK0ddUqDN/WOSkthYSKSbG7Ghawtz4+XWiF03I2exuuEOIyaAmWGV9cfjbqXC
8fxEq5I0K/YsO+tkeehGamg9/0hjJ2XgWQEXtcANtL5rShqSbTdbub2wfDJksuq9
x5aJaQ/LpZswb2iaUpej1e51nM3DAQzuaAcZE6SLihatahC8PQ5UwPmRDCb0iH6T
wMk4px+rClXeQ+a67Fc8VLUycKcTjXAwSh7KzEticn6cq0nzQz/L1dnW/1tWHNuV
L9R7ty/7Ek/ABNd7Qk19zmVuwn3qSb/10facFu1bLAdq9/2PUWxKWTVpRqwUZgeM
EgHzSfWjCTnldicdabvJbRosUQzLYZNdTtLx5yGHAKRynBk2Fdr5HFJw05BrJs+6
ilPAQ7tMo73m4qSEXRDFhiAGFJjI7lkLAQOY+VLNMd2INCNhANRfLt/6AunnqIU0
t1N41UEga0FG2OSK1dWpLATvUdn8ub9SZ9cYIm7hiUeacwiLCCKPORMrxAKyt2Em
gKYNWaYMbzPzJYRKYfPwvzNC3Lup7tR7mTQOOJ4klwe55cvvWGdXsYigHPKsvgLb
T23nchMF1PiJRrg14S9Ya4upwwfebApuVbeSQDN/Tf6YfZFDCuxoXtpmwVB6Im6c
bHHyNhglUR3cc66wYuRvFwAArWBdmxgewU6RG8trly/abXg5YCsIuXcmgXttevAt
b00qFfUX5hCny1V/8bzG8Q+Mq/BfK2W9+S1V57nmAGUEStRXGInHPCgrxcc9xMUX
Yg4a3/nOT50RIpqfUn0d/ytefV2SYedYGAPI+NnajTBkqtKrjzQvA5Z3RkLpockM
4DEZJbMf/3ogL8D1tWqD0OoWLQ18S08k1BrUn8abnzwYXkB61pycWfN4p4pUO7OK
iENM8CT3n7/CzLgX/nrz3wYZPnvUtC1ZpA2Y9polASdFpfwpcJLQlyvn1HiiKgHp
oGra4gkyQyE6GrO51Rvgd2rK1L7xXi7aAXDaUz+XgG2t8IflrQWxcwqviWN1xBat
SMJ8ozb3FeMLDEq2RI1VzwlNsuxqIedz5MM9lWVOdP3R5wd9cAHdip4ILvKY0Oc2
9wyTgsaZlDql875uBgMp0Y0S7kk9nRZlvblxYVsiNk6Plmz5wXgseLu/emrrAlFH
Lr9LT7WJ3azAC5VgpoVYe/FDFkhuEO89ChBOVM+ZIJjF0v5LhOqSFN8tCKKEt7i1
91DUBruGPOvZ+oHM6oBVl/xNcXcrN0uEYtbnChaaP63QSal8iTRrhJ67bTerEqDJ
IyvsNAg9Jbj1kCnF96zIAHYOPDEYvMbDCn4Zy+VoKXr2eDAHqUERrjvPzHjpte1f
AGDZm/Y5KEh1Tafxn29knO1j0gpWaPixpw/VJJyg2WtFUAL0NKhrtyukIaJyXMEi
LKfOZLv0Q5/qhCxRpgEXYKKPTje8hb8c2yvEhvprGDFEpYsguMo8kiQNmeC9QNpP
bq1ib8V2K/midGM1cyPiSv/Pvwe+BbrTmhWRAXAUYgl7hjYbh5kF/nfKB2f57rWc
15aFSR39hYdjI7+cMOEj9nOBenVWqzJwAXlhR0QEeAPNm5Jnk/VmWNr9wcEVVcq4
8/qMTYztvjBCZ4SybMQkO1igvdWmtci9l36LZL/5j6cjnzli0btA2+mKPU9hJf9b
CHSoBj59Yh1WgsEtSsNXBX6mQkLYduUKKo7cR5/IFASLKSnt8ktVMGUEZlEMDFE5
+AJK+Er+UA083DBNQ09EcB+eVX2N6hf+tar1HiNUh3mDdvREdjno2NyYOdUWRsBG
R5WAgyQNvvCh+cLWubnvMqbGvBdSMGVKcL3C+6v/MQzUttzU/vrXMYNjNe36OoDN
PdzKGJSqrvZVpkd6NUubsYiHe/HDeeLPNHCnIrCrNSA+/HFB2L6K+uA35k3DHZB4
VdsZhuzN6vsc6Sx5z2gUsHlsNfqQp11z5K5remEjrJkTpvqZDOgqzhb1+U4lw1c2
XUnM3crIwVtUM90rbEcdbAil0x9TQLwRHInl2eygLFw1cKPldWjCa5MV9w74R+wL
cRukqD62nG1ljkSDMbyMNbt/E2sU2+2wHGvmguEYcrEftJZ4tvabZfn7Et9211aQ
5Q0WbRmYL5r3lSbRprSMGJKIxXS36xhsDyt9EUAhFGFXe+Hhlfw/gUecvZZRmROb
5tK7EI1HerLBdh2CFK1f40D2LLdU93Nl5sbbmgdIc2ck7yIBKMpxKBwTjbQf3CKc
ScDyJlKTwC1BWbLBpKSDiFUcSuwJcw6INE9MB/UvJI19DTsOM29QiTX4XlsZ3NSo
jik1n/hNwFdU8r7wojU2kZ55q1n/vV4mglfCAwUb/Nh1VBY7g+nELGDwSBvZSCnY
t+W7Z6p0wwfEX85fKezvDlGKMbRIKjEVZGiV2x8ihN/Pa2pERHqV0pRV6ctAzlT1
0CdqcNfaUGVm8iyHnQ8fFOCGIZc8R+9+qviyX7pdHTDLQyOOO4VBpA8DFfink79Z
XgklFKHfe3dNByKapqVdZhJTuGKfI4V70gYXPQYyIn3CGSEhEX/fp4DgFFLBDa58
Ij/Fb80ukMSgv2tvKnMTX6pPrjNj2c6/AaZ+RF/hZkVYazqyGn9HkZvPCiaKEcqr
MWsy0GKwL+T6YzxivIOJ40EGoEaHfg9QWHn6+OnMkD8b0KjVAlPKDcKxRTKmYZYg
taV0PUAM9VKP0O8DV0ykYWTWLAl4KSIafVKBQ+vmLEn89I1xC53tKFl2tRDclf6A
bDNmRipyfZmDXBY+hedhMRSj1OPOPgPgi7c1ndl1Z/0u/s8u778DTMGX/MX2Yhx8
EpIxgogtPGsVCuZF6r8+uZ2gISZbEHuWaXQe+ogiYu/Z/mkF5BD8jQvo7G4ldrV/
JbJAYXjfuB0QRCmYh0rDjt/EZIOz3DfFNnXzH/tRaJ0=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
g3kcNRp+PC+XG/jRVs+YSjAXn/rYg/eDZ11J4ptW7qYVu3WCsI5SeSECW6NSh7jo
9y2uRL6/VQ0d6U5IAehgjRHyagufkjJD5hO74OnqsIeABLJd5IMAtstvQ8336qoE
mgE2BQhu/pBH7a6/am4uKeCegP/wsBAQn6KpajrYLtcw4NoCAMUhHtGCsSenvxNM
DJ4NxpO8mmhYjRY5M8PgH9oG/H/x56gMHpDj+nIdQYeS4rzysiGZVYsGs3fJ9b7M
HlRumwR5U/WkfRz8Wzzf6kpDWVcno2aGLTLJrRUJwQdOC8fKs1rvVchpakmVQmhH
+i5+ecUMgIIDJpLlKiM4qA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2384 )
`pragma protect data_block
q/ABJICxa5GRn5pG+OGrJb07L0mCufN/+tTv750Ret8uwBckb/guIgW/oBuiuUrj
0v3HsVNM1neFrCquIifCkvexCfbOftMjZiLwHoIdHMN2MsgVEOAJjQiXHDpHRC+E
id9i45efahHfinOkkh9T9X3K3tOy1kGBvDX2+SP9I/3wm9pAjqhv697jDL3s6gMM
xlMZ9qk5ea8mrOVOgpsABAkbcZ1+7ZbtjAjK/jKh4sF54fWFUgn+xmAQ0o36h4e+
VVwyS0eGt8m41Ev2iSVdMKXQ7Xs1nDLOqFLI5esHFeAhYGZZhcqzwBHu8cCLCyWi
zJhi2pOSVkASeuIBtrZJxO14UYng63kSmnWoRy83JPR5Q13fYjW3o26a1RkkXX8B
7WEDqg3I8KCNMCzD1iFVoO3SwME5RbdncvASlaHGgcZ03kxV8H31zUcjU3Kp8m9L
fBkCTRNg+u/ReT4l6OigNsGElHklHlA1WB0BQi7AqifUipL7M/HumRWVvVI4pf7a
/Q/JSooVCdyVJoOameo33cMIzAHI6kGrgbUX02rHkv0ZMrp4hanifkMfyHAyef34
YFohTEhTSFOsb+lFxTnbkAJWnUGMDhB+04m+sRO0tzDQVPfZcrPNMml4LjW2DObL
riHwllWaVt5V+9JPEhT45zX4wErOsDx2XUWiphHNCw7EwKJC28bnXpVJPOq5ZLr/
uvkHHR7VNRPaoZJDNaHrxVBZ+Bpqn+er7RXJs82U2WPlINH3OKUGwpMeHVcLmqLF
FsTlwvmiXKUHHkNdyWHQ9QCTAnX5DcRMj6RUeF2hfh0GCeibLQ4c3W88VB/7I9nx
7I4Q4dyIzztFOXmFpVEupOlNhrJXbnSvOHJpUvHPZVHN0nveRoBaRiWv9tFVhZ5k
L4Z7i1Ne3BE50XZnJoYMsYymo8vSJvbzwRF3tCpgF6HcL1gk7XfHKyTVD6H0HDgf
LR3LpquXmKZt0DQwpFtz5ymro3MIzjulvJ43/BW9OmCWM8Ezn/IvVBukt+63mJGx
zgvJRU5ho5yaOBIbTEWHIpSVchvBLz+050BJpA/hPmtfgLWLFznNUkSUsgc2K/gj
VJ8BMlCWVxhBHFOl93TrCB/miaVnntSXWZgLWam+MSkXBnGgBT7tPVp3Kyx/we+I
Q60LBh5kUMFB/HhQ7UYG1DG60cLLEWNKWlQlXcZ/Gys0/hOt53P5kfK8VggNFFAz
CRJTwh+01fUc2xKYjDM+tvXnQCsDKtFZwAxxn6HaTE0+LPs+ygXV0pCsPSNhRBz1
5uZq99pjTmCmvCEtNwvRt9StsLuRYOomwtiTRS12Gg7E4yjisUd6wuiRenv3Cktf
axG78Z3e0ROYw5zBGqi3pjk0hIPIGGgR71XKKXw9ai+MQ5zBdCGrsUWFnrOiT50Q
XvNhr6TBY42xs55jPyuqAiq8zRdwpEIqTi4awnoLtIAnciYcr8s1l0QmP4IFr1PX
MDKosPFeQenQ7ZLYKIajVInfLLAfPTOmMk2Obl01Oop2/8Hp/gXfFVNFU0vfSGx9
TenZguS9npfo4TtLOl22V/i8JgB/NeM6JM8EnBayNlQAu/924WMJcmDp7ss4zKG5
udNwJ2p6vLO62PSp2v3F+UWpdFtbmA0GB5QUXJo7Du1fJLi3q6g4xcyWCjI8QvO6
yaR+3W4KovvXIax2HEmTIvhSJ3KkxGtcNQI5/Ft/dnw/LT90K/W42T/016IJDCis
7iS8B9AAYJPiwYNtE6KCLj84JZrwvUH3cJ+zCUZ64acNqWjPhpi+Uciok0UsST1a
VL2P2emq43R3vP5NWd0zhqto48zXDKWI6DBQ4zPO/EdzklzGV71C0RLQAuMPnfl2
uu1EYco6wWZaAP+rRoLQWutuPbklDbbyGhZRMhEO6Di5m0jIHpwGZKTS5Bdlgl0D
BHq5GBZCg1tkiS7R1GT1jZ5NtOumu8QvoS8AHWlsxkJ+PrLm6VCjY0mViRRAdaJI
shYJt0mmoSfaknemMhmqlNwI9XmYY3tKHNkXYLPRXlBVgXSqLuEMvDyQu7XYkQsu
3rsnO9HZwXJGQMZpczwb5d9R+WuqfAZzH5IM2bU4ADJAwUA2VqSktX6J9CtzpYCk
oH2eb+HX3RS30LeoDrgKGcfSLcODvJ7B087K8/IFdwbrGKVCc+WfRTTXekhS8tZV
CeHIV5m7U8U7qhr6mz6gOSNaDOFP93XhqmNwJ4s5egnmMttXDkrZz2mXXDDkGnw6
18YLJPRl21ogJROkESp193eNg9bYzlBEWyrtM1GDB0JmiiQuITvL7Bu1ZvvDtnPu
WlBrUfa6UZ65v7jlY8sgXDaAMuuBSXdCL4MxCjE8qvkbUHd7xQq4H0KbJggzqqqX
Eb/ByrNEKjuIXQj2rlUJ7Gb+bz7AbNe8a62CngGJYu4wDUziFQAy605MOrSyH/XG
3aYreXWIo12R2/2lTIcYe9Nt1vRCRVzylsfIr7d/tL7/AGb7qRQhC4/svVWBpkrL
SD3Q7nRIPdD4AnTJYZMJ2XeWseKZpEq/rldQmG8r/Mg6L/sqP0p3AB5WJMIK9mU6
GCCjnQHt1MghNrhvqJLYczg50Dc0Cz+NSux57Sx/rvF44aJXuJEWxcb+rfBu4zKX
rCjCjrZE0rgdB1CF0jK7Ua0X615yl85IQAigL0LDaXAFUxqFU4vJIaW8DKqOdJXM
RG8q6+l/ZgmQOQx2+cum//zMJ0yFlAgLeZnFBUVFV2cVVNa8vbEgIyylSlufh20P
EAzlKl13v/Ge+Lp68vYCXZ4qeJ86hJ6uHI00dNXJzunZNOefunzczgEjHc07miac
PNoN1O6ZWficCIw/xSstKOnCSw3zseiM31B2QaDDZHxHTVnltHEIAoIaEVfp10ad
AZhccboQzlI81xGPBiINO3u0fE1koIOKqFdNbQvIyiORf030Ot/T4KRtuQ513OMt
YrHwVWcwOgZNzawR3NgU6cH/nHyOXCMHLbVxcMccbhyIPEsOM/kFhWOL5AafijjA
XzCBjZc3v0XH6zF8ERIr0zyq0qhvaDvzpi1+VoGJf6wpbcJ+sBDariCJkj98OZl0
rvxl2gHdMGHa8vlQFEmdoB82eFZ2jPSZoi/XC1oMLLtu9x/wYCpnNL2wMsxTQbKM
bYTxSaqJ0T7b/oOpr2XilUNg784sv781h5lO1mKavf8=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fNYNC2bISgVZeEf933FISqxPhQPvpGhwHAyqG+NXU2bLqFv7PzqFggfV9APfA4U6
ablIPnWTJBm8ZsnXpn/ty4Rz64Q5l9yLNxPL1/Tb5Tu8kDKcO1Q/WQLiPG8I0SyM
FhdMpZ1u/OGQGE0iOLj2ODd8DswloFAA7nJmyD6LUeo6rpykqpouJES/HV9RyyMl
MzQwTtFv6FLYUSef/iWjRz+PAqSUN75nQU2sHDW921vp6FMuUZfXvAlG2qulfDfp
w24aXiiPY2zox/REcSjJWMUpiGO1mpWeJAQesG++EE10hqjYQaE4ozjjk+twygcB
sD9GRkZh2t8/AhOFAUIH3g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6640 )
`pragma protect data_block
2SVN0eIP3IG2Sj9JwKMUKNFzEgqc/vIpyt3rYhAYquqvTrgH5IdQP4aZYpWLTNK5
8oXngq28uLKRgP8NwMmFB9hxYLtqBJjZmGvsr7jnT+Wzb+CJR6uBGNnPaXVUBEkx
XDTvZfd/uBeEVmUElQjJ78kNE42UuOcR8ATRiND4iLDm91QCDujwV0UuQX3Kwjbi
Ezq7hJGJlvQzzzGGEJV4rTC61IjVRfFq5pMTv1hNsGJ/IIABqvMrUVDZ5f4rXBhr
3mLd5n6f531/3Z+PBLgKCxIC5Vd9XLThwzWRUEgdEKQDCf69dapgB0bR3IUgr+K2
uwr9i9EsEKJfdy4fT01toeYRUwQKXEkUEYUKqYKZAXeyo7OwkFof3Xt6tNGh4Sz7
JDhqxXiDpaIayGY7gDps2FLSU2VeU+VIW+sIJn4H/yNCnFDjcrCGxOZH+mkVcZ/8
USaJctu5J1qy6cs5Ct8b0gk/hwERX6KBTi/kf6vLhcsSdvB64RCboFuhkJhE746t
yOPuhu3XBEx9pem8SpRo1QI+UpiprOKbQgc3OexLnzSIN5d73QQwSF/u3kWbzBI3
ETCiG+I6w2cSaSEqyhqgQ4I9iLd3625V/m/6TJs0h/5PQjzSljGUi1dkN3nyi+yf
90boZqo81VeCBgMI+QPrjYxRg3mnVl9kpd+UuEUwlsK32lXwz4bZG4lrb+LQ4h/f
J7w22STmWzWZw3KCE7uu67D7VNMW42JbVHaZ1fOEiSz2JEXG5gJdMSoRjkwEsJPE
/8qeKqwnTvctw44SLtFOYr7egw87+qwqLEFZipqjGSpwMyQtrsAqstTsYrlqej2x
wWj4NGWl9UqpnyRLCRwGAKqSgeYDyXrgvslD5MvW/lOIY7XrgGK7ZojaBklZNkIK
PgjUnB6ZAq0KFR62c5LuglXTQ7E/mWccEbBk+ozSqOhmcLAYOLCKvIGqww81xGzv
sU21c1qYCHTHkQRuqj9Tx0qpP/kyIBL1smfmrT6Zu2Vb5C2VNbWXZ/V00shy2xdk
NGxdo/lmhfbtDm0FfH+MtSQtF+PW0Ms9DIWUpuIArMRp0XLwj6Kf/HV3aXJljAxM
A4+kg6gems00Sl1SEjg/ySVDtOOYYqS6bHI5mCPPV7mqutsixu6K7PREwOorv0ji
4tCJufFwfvL0zMPA1CbhgehbPoNuzt72tCdXal+o30ElsuG1Dr8RBJBwg88Ix5xd
O3nlLUw4PFr9J/bzD+q8aCyHClOtSlYpzoZBUCWdeoo1cjSgdvNvytr8BRbuC1/b
RqQ58xVwpfdAZXdJoxbKdZmwZWY5PCRyammryRJQwy6PHiojv6rIrDzua7HzcIEQ
BT9tq+M5tfCkc7BIq0Tl8nTbYYlPc0qpk0i5/Cv2WRUDPQtxYh9hg1b4qOBk8sWw
8OXKRCaHFmN1sNXleLfu+C7vi0UZ4H8XNO7Fwq4U+UBREwp9796o5amYMOg0yAuM
FwABlrCd54Hk40fXmSKRgSzDOKqi0YBkeciG/Tzj1KU/eLF9mEFchpJ3rCZoU26I
TvpJRf0zREogTdOt2NO8upCsklkk9E8aQNJiwqQkUpp3qUSLzvDyMChlFxrtfvtY
F1JSepdYUPWWL90GnENObXz/fFpseJWZgrkLu+wJJC84+3PS7DiYiGgAH4HNe6g0
e0TyrICEKsFR1ftf5NtOTflLaYBzK6pbOXfAHDcPAZeHZafRdrxtFYg6MjGhVSO4
oh6puhXwgLT2wCrNdqe6VdRDvx7l7G1ZOvt/tAeBDEsTEIgo+qhBsZO0S1nOr7ko
wCyNsWBPNsGk8Lv3I25864nrFfqDWk7vM3GoOZhxoMY11MupJSXftyaz0gOcoYcu
3XCNjgGSkw5CxiFzCWAJoMP8ZmdYxmwR01IU2R3BDeamZkiQlN+dV8u7n40VTBLE
gnbp5Gi6ICY5My734zinq1GLEG3Wuq6PtxMy6+FxCn7kh7UMxK1Kna9R5C3lJO5o
806DkQot4jo8NsMJ3fDzYxuLc8xr2bOIiYz44r/e2LpqJO80JP26kz7gZSdFjuvw
6/lUvLKmhH4KFTX4qS+q1iiv3LkuuK185y+i+k1p/2I2rWfODc8fSL3iKEULKR4F
SVFHfh2IDuwQK6L2ERFnLhWbpiuDKATvWV9Og/C5ziroV1zqczlhXeg8QGpd/alx
tAToR2qK9hDNmeF9B7nn0H/GkLArndxa3jRu7f+S7n6yo1ba3PndqYafJVOpmOlg
EtASUfen/EBUWdYsOvXmChDSclzEeOndupnzkdbABhKs0JE/c5guQGH8gqnrKO7e
Zz1RkVg11Rj3g20zNxb2f/ZJh5IxhG5zq0UCn4ZAFk0pBw486KlWNojEqqClaCfh
PhXTF1StEdnThgO/YnZfOH366ezWS+2m7mcD/uG10h0d77fxdDEvRsMPizz3yOos
lAx/vMnFmFNajneIpmBTrOD87QC4y/xwebSFI9skyrx6L2GXk5JaduUethZoD/NS
5SLgFIy0X1eo7QAJLYycVOo3ufosOELOONYy3J1oVRnptySl0iijpskiEFYLVnn9
p8WqDhX30WZWVprHiESn5CyDkgA0lVIjfRwfkdz2v7gcfIfI0bJsSLHOks70SPLn
MChABw36nXPS5gCucGA1/p1j/PAU0g/SZeLRG+wzLoIM/GqAM2hCd18UkhiO3Q2d
fIbDoY0eN/dOoic8fCgF2J1EW2B+t+sMw1lzCfCfOK8RSyoXiT+SKViWOAYir3Oj
KKN+JqFpgV2nwsFXN1bHDuxIA8r2Fz/2WHmMMsVlexaBOGRBoJ/FX3JA1syEaYtc
3EdjsaQqK5SxOx9yIAnIMNiKY0KYyUpqZVsVV1W5f/uS3lPPQ3kjPIHxukWpXjx0
mekmaCyU5iMGhAN3m1oR6Bu74BXAhdB4hGmk3Hh/4Su3Ma+sZRk65BRSm04pUIyG
Iy+CyqmmRPDvQnOSo7E/SPY7QMTkJv9MESJghkk7nFFNpfMg9ziPjUiMoD7xMEKy
s8NZke4Q3wBFziOUWMoQctPuj/1raFzbiVojYW8jjIi8+Phb/hzRQXbiiXrD3SpB
jYnTneYsaA2f2El3qKEQOUJfMqbKvZzpB4jrje20EuH4VzB9LHMUaWhc8cYnLHrp
g+cm44jvRaQNKAtec2uUbho/kEe5nzKpQzM4XKa+nvDg+vp3sIc2SE1RIAzOUyNv
IgbYc6W29kyGBc+oqNg6I2XpUP449pgo5WytPCOidmkfVddaQJ4EhXpcQFz+VS09
zRu9CH5G/XtB3bew618Dj07lk/g6uiLdt6xnKdapMb/l2F+zKUbFa9xAXXS+pjfh
1eisUmtSiHK3Bq4OvFL2SIzIISNdqh4Jq4Oy+IblxfNI+JdMYrRBZyla7pev0ulA
ksHFH+xU6lcXk03p0Tt+Ouu2p+9txNs4vAd1dhBi8dGuxXH9nx5JqbN5BbI4rzdX
BVUNeR8/F+Lmtomg00QNvxbxG5jwG7QeNOYarrcPDzWnI1UHWKelnyzlhNTw2B54
40jEycGKTQhZrtn5Suyt0xumNAJzRuOlHFW/zMl7jf7Gba/Ict2cPzcNN9pQDSkS
DAjCbeh6CORLpqSyjlHSun00LhFsW4LvC4UxluDolcMpw0seqC9ip1+ZWicZ0qJa
6FbiHnq7TPPwglNAkT0e48/XhOIrfwPziEAgLr9UNwyt+IqnNS3G5uUys/vxT5TZ
O2f5ZrYEsl9IfpALvcu/0JBGII5nW/fph5nwJFWyW++giWC2gSLgb17yD9kvre4+
5btN2dJNV7VOy5KB1LcOUqwC/qC6cHL0Eb9DlSE1Xrh/OM8EaJYPA6Adym+OA3+n
GN+Q+lHd81j8XfEljZauARpsKWYs1HqIB4fljN3WFW57YzD5tNr0PV6kS+xhS1BC
VPjeR+5Qr0N+vvrN8FL42yM5/lObckoskbxC+D9w3j57N1JYHRfubeEYb+3rxlZh
H2OcG6dELUc7tA/eZGXEXgXRxoiY067Xv2jBKd1fAiw3ZFVeiTCUHL5ojN1GS9Zb
KeG4nq3LBGjp07VHHHlBsEmSnUeq3h8C1ouY88eetuVahekk/S/B/cZ2D7EBU8gd
6LdxMpc1aS5XnfOWlNf5pCcX94n4V87S3pVUMmGeiXihDYlDl1VthEnq79xHGW3w
FUE+5uuoz51HIXz658/pSB37zBd0RzkIffkYthoUJz7oGwsAgJGotw4BSGNUAuj1
lHMgaZbDX8sTZinLADZxSP/LvrcGzeQtvoaFa1QbF7ycga8PTdDmwrMykg+b6Gyr
wTgM/U3u0HXSeyxIrnJoYMXwiLveiqnhj+lgy1qkVgF8B0jSZSTw4xBiNbhZ6vlE
i18ohCmA4tZ6J1hVULogXOrksy7mOwU6jkzaJXdG0I2uVXtZhRm/3MKsqwqA/BV1
BZSWy3S7hmfZ63/8pkVtQzTRRWuc51Fymy8G6eSWpXItqq/08m/6CU1cpOYp0e4P
i/sTFsKykExRRaERCVLrKOM/PhZS1voRPhTsntS5drGET3wiEFygbtpBhe/cm3V+
M07VdfPNEIvdPPKmwGgZxCMUreaHca74pDdMY4S7mrOuLX/UC/ytb2w7skWczFza
0FFUIAPDhInBTPpZ+jASmK/C/dG0B4q/wVo/cdRFM1L04QJvmfTv4sM8+/P9LwP5
ugiQ+Pch7EGtSREGecHdKtszDT70+QptFTKkotlK+L/7B4puBSKhAs6ZlQivXbdn
KnBdUAsUyzr11WCROFU1wPe8l7Q+0pobOH7fW+F1lEZCtM1urr9BgGCnwlHo8+Pg
QZasNv+D9wR5NiGtKPrSyAKLnpkZwzV6MlmFz+uixMMNYyS8kz7Gjl5Y1cWUpZc8
OGfSxMT4+ovUxlyH0kVDMEuCh7QliK46f95Dx5NgP+lmRBZnA+koqrNvnpOoIPE5
eV+IXsSKuwW5XMBgWqzV9qIdSl2AALBsPiCNocs/WvO3lSXmLmtxJ/vJPLTx86Cc
vGkckTJfyRXiss/HoLPEGMGpzZTIZqUSrtfiZxQ2uzLakuVW2ot1d/QjxqTaQeil
6uMsGPRvbZPQ5+51DXczV8t/9I41wNOmlTvyKtvataTxC5oO36lFlzTpHDWruMvu
l7WaUl12VtxSt9lRhvKRuoDscBC4Nqi5Oi0pKMRPTA+mwB4ZZNX47RDeURI5L3Ft
TULf/BfaRL+iYKrDNZVNCVDtTVRKWfR2k7d38v44jL4xSPh81vNEIUh7Tb+ESxUD
jpF5RZ8kh0Y+0VZo2t1HFAJp5CDVthU+b7XPE9lTlVvrKI/3x5U+eDEbQ822o0q+
cy3xKQ4tfPIlev+Wn56BltAjDJLjZK5eKuPan8kc84DxWz/R9a9y9QiYkxFEDUmD
XP5SuGzGUINeA5pmsi7fFnyweDvoUeXkm04luuL5nS6acavuFci5SKJgHp6nRT/b
Ct/q1Ayq4YmrIxzOnjeI++lAVjiHv8ojzuOVZ9LG3pXuB8ZBJlF0MSGLVRLlVKdx
PlvuR4anu/mFz/ETTSTuTcFvLA/fY8ZIEatxqVwWh/aHar/JhcQ7CAaPkP6h29gJ
M+hzdFbH90Azdd8WGt3kjJLNy5GSO7Ro6peJQ7slz8KgivLCFDxsttTQugEF0qbl
ym7XmAHiHbjxXWBIhpldXF3BqF+7jSoRhZgO7IZPxYHeAuONRmkVgpuJVNZ2AWJ8
A8X99cy2MivBofLj5cojYhAxv3SlwPNqgKO+WIPa4qMPiDW8O8CQVIW+GqH35vtQ
EcReixNO4/5xpe7h8cUaeS3weW1wvaNuWjGIoEnq3YYrqzMbZpbWjVWKLAqLStkR
YThp4jqc0AjhvjRiltZs1zvDbhEBUKO547R3Ibx58suDlh0M+X0pM8SLT6PKnB1a
efHQm2FX5guCRviG205vApvKfsJEFinQCpghM6ahLrPgq25wuWEEyBPBV8SlFLcW
/j/UZhYF3EyRYY25kQJSgFUTkBcQMTsRlTMTEN/nSRUVOY7N0p7ln6BYQ8T/Z0AB
neAeJh8fKXXWkdrDTtAMB02r4kSSfSVENLylkF8ok1tQ54p1y/UOLrbcceUKyBLl
jrBEf2QmeUWr41HN0kfaCrjkhNFEEMISV3e8jAgxGDgZ3RLJPcRdolky6c1wClzD
dXo1jtzRWQAaC9k49CDx0C4vy8RhCmowjylnwXg8XhMp4m+BsFH+xp7dSUXKwMyV
YWVzHvxXmu81yBRPRPm7XRJW6kzorZDPyNSDCu0WbCRf38zxqueQX58uU7q1Zwpw
eqmwsZfV2QS5STQqLmFHCMTJ3zMoaTqKQvN7EpW9DX/HdU3t1ZCEYfcDZkBL54nK
fye5KGAP3PT52/Ri58/s/J4fmQAAiGuc8ReAceYkTe+XXlD9p9uVZKXiZ+1QyW6z
qhs6tSjvOpKK8JmsJIffKwFJE59e5NtXKW7JR/eX969MAr/wLccFUeXW8YD9KJ/k
+eFeX0WWJw7mojf1SLNmF4hYlT2H+Q/TS+PV6/k/5VjR/KuHbG8BvjROHXg8ScjE
o5z4FvM5xHoKu75HyX6qdpx7noTt9PPzHhqhTgvrGCo+/VkXdeE4/LYsqJJdJr/t
xPwdkSD5AhUaWtvd0Onc91qsC13OVpxUZxRKLWcZ0xRCDht1kKxSv0e4Nzxgs2ox
8mjLtM09n24z2DmvDEWNgPuZfJx/X/C/g5seNg+5t9caK9MadCbz17hnmUcpiJGA
YSyczaBIxS18rDpUCeMsLK9awiWTGxutePU9cABIvqAAr2z1coLC8j+LmYBL82ZP
yEgfdjha/QHCoJFTc4nB09PDbkU87xGuEryMNMSfvf5oROQmgYjGWag1zoYeqgMc
Nff3+LBPNBzd89Ob6rP1fWFJTBm4l3nGMYuD69I84DKpSBQsH7Edj4pxA8MRMVLz
dMSUZpu4ljYDyB1oTCyJdY/D3XlzR0dB8Ki/fD5RXJoNTco4p/ISUVav1Z29LHpk
c9AxqvIk4xKXkORaqln9Ss1IoZjctWAAgwxV+Vb8kBEu0tBFD6uL21IdzCrX1sGz
qdORRIxRPWk0hGNE/ZG3SrIIeWTXq5GT9c+ru4ujIR3MUZGYRHS8MdzEaA/p9imn
O8eJUGWoevGvZj0bwW2/oMt8ANWRIusapfwI5MXbCGG9o27TaHXCkDhyyS5e/6Gy
35WH4OSNM9I+cPkFwzSEGFoZpkI09FERwOyH+PAI6j4gVghqhai9IOJxldKmO4jw
zB/ihpZ/UE84TNZbt92C/dLem6Gt9zWWi061/agzGsUrluHqf5KL7bEwOISXMTXK
TK75i341+qdjOMDpJouHNZ8a/WsjMYzr1y0E3YJ1EkI8bUu6Uk3yQgg0R6zMWWMd
qxrYkpF3fbsnuxzFQkQnjelN92kvg/NdphYp2dc4PQZZtYVvKnyceDKdM9AwI5oR
1xwoX3armModHKZu6A5PSxZp9AqCkvs/7kqu92CQ3LTDR3IVVl3zlNuiTcENLAJ0
NCJgpP2HQ3/omFY80lM9Y94JNv+S2Y2IwnQnk1bRVSLyE2Hc2kdsqaDecAlRp1jd
5MGYoH9YwzYYl97R58uKlqRwnq/iFZrTKeo7X61qFSAiHFOQgvVvd7Hols/QnMCf
Ynxf1EpfCGQUrBj8/W8fw/gamNlk77QxJXVrb2GXYFT9G7HO34Yxy1DtGLjWaoX5
bSSjc8HHWq9VBl0No5rkSy4ctXWXP3sXh3N+x5Z0d6k6aGlqDORCVpdWleFTsRu6
PnpCkSVafX+K7p8K+EsD2baDK8Y2LhjwMArN55fqUj5nD1YG4lSJG8Jyp8YfX188
RDjmPi1AeFRaDwB8qkM+4TbzZqYG5RKaqebFUQEsCgNkwt9XvwS7L9Zmp6mAU9/l
06CS4yOC0PjPgN8yD6Dnnsd6ZEDLSajgcNWuZy+I6EcSx2w5Zc1TTD9WzW1vx7hQ
CKaN+BraFxX6+r8wC2PVeYY4VIycyB/BA6H/6RADC/TfqyrvgG5T+789F2VmQDmP
cJ9LsZYdpLllusHuUw6clHwcArFa0ybtmGX7RzFQCQGT2do9pmDVtqTLub7Q5GlC
0inMj1qimUd2OkWoWenS2FVnsbfPXf+wDm/Xj6IWLmjbXLIVUFhsajro3JOHL2Og
a8OYto8KxTNv5Z7jfydKIoFukob8XkJ1wKpMtQ7de4fo4QyWR2ZvVGDTka2pYEMP
wD96e/Xly2AyXCje/D6vtt1p0qM43u9WLw48RRhdSt/dRqg79jl4iv2dXad+HHKo
8JG9EpG6POdPoZZ75Za70s7XM7T7MDSTQ7tLg/azhGQ5zVilioz1xOlntmSL5OHs
h/KJlstPxPOFA6+oVW0hxQK35cRpo28Vzz/Uw9Tb7pfJTEtcTatOOjgBtUBhRrIt
d4Rv8VGgzsk0fPNyUoGO7QcpQKNIkY0mKcscxWLgl9v3Kdev6gHIWA/Ldn4Dl/LN
g3RFw3uC3mGTwCqS/7nRkJC5P+TKZr2f0w/CyaEpmcujhl9gOP3Kkjw3S60ZP5I7
g2rhLcJ8AyPoKmXL02djoCqp0wYLiAHj0aNhzfVuG7tNItuaAOjqm/l3RSLvuWq7
ylctkLXRRYzh9+IjNpUzIkJ3bVyPMoKLIYeTOgRffiW+BsUdArhSxwsqVCxwoc/8
UTembt19P/rXYNBo06R0kcHYPo8IedmDqtEvj0erFojjLpTpUWm0nkzCSwrb0H4V
VpCTY6mEUpghSGDtSjBr3vOUPz1MtLcBA75Knokv61OEZn4kIFD5QgqQxcqot3aw
ypOZ4b8je11X/pcKmi6cX5WHg2Wkj/qGVe/CS1hrb6CBhdm332Kqs6zCqd8C+hL3
iAUYNk6Qc6Csi16nMqEE5A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
A4Qc4siChBPK22lgANnOxOEhOfl0WqfFT3J1fNzUcrVIio+uLTCTO1CHCIN0+RjL
YnbNA7xBWDcBiRcyDNvYW2oTmU0fUYO1S9K20oS841Vi1s3dbs8s4dE6Bkew0XY6
SnFpLL0SlLyVo6iqjmnIBZhkERENsI9Le+mWuI/mLukUrcUsVIqj251DXrI0yTJm
lD3NZk2Kup1E/d36gMSxUDk33XopFzHqj0xkHTdaI+VW88QB+3XDN1UqZ0qwUtz6
WW2fpYwjKsh37JWMHQ3BEwHHl5LVrVzLVWde0zhc5U406P5n3t6+KBguneHV4qxz
xLY4z5mWwrdNaWjiUpERiA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4960 )
`pragma protect data_block
haplKkIDOvv7eAnO0jpuVTO8Q7OSSkzbrSCVoYnJsgPcME2BeilpmjpQGctxFeaH
7sh3MVhA4iLuBCR0zymYeaGqrJomb4nKHFVcMFCmxft/ekNI1wW+fhCV9T55OyzW
3T34k+HdDRcyY5fpuObYL+HP6xWmR10lcy/XIIfVJfXjli9AYEV6DCyUv2qFG9aK
lIW0VbLz45t3k6FqJsJndwdqhcjt5P5lvB5DFk3h/xWmjJ90FzqO2dhb5a4Uh2my
wC00hynbC55UVHLNAR03drQCXy3D2FOEnRCOGs2cMWgEMPFeWQvBqW6Vji0sFoi0
07aVJ8TU3z22ypwY4h++AxsEC/6rywf6Q1919m4WQYDNxIv/M8AaiFf3c42GX8lm
z1z5cIqbusxD3g6ZQU8zBmA1ll4EUfL0E5K2I7nqhf50Ixn3PVr7qcDHQsZpelhT
/dyp8SxJ+aRDHlDnXcEKVnftF8vwHLweTwSL/VaEtnKMzplMXaVlPtHJHu8BGz/7
Oodi1vsnWfp4MMCia8b/1W79S9HOVskCg2XqeN6RoU4ynNouLwGUaeC3m/8qaLJ6
ETMYLkimy2tmSjbKk2PFTJmf0v3NEcfb5GFTNtqP1ogDFRsAtpkiqeH9Sg1doC8z
ICONMFstLa5DXISrDQR1jQTs/AqBShTUflAsnTKNJdVn+58G636JnX0dJvwCI4Ef
fIB4tWT5cyEO7+2tSJ5ZfsDDfuCIJ42WU+ySX3q6jYab+m/NU2sG21RmJ4jU3091
pPLIAj9NSqVZRhFctEK4Ave/UA4pa72CIIUZfZOK0tIQar17cJKWmAPQD04XbGty
7XcJkKlN41NVYXOp7Gb834Jo8QlMVr05/pGHRoBDwPjcB8KLodAYVeO/dWyw2xtu
8I+T6R6DfHhARtcsjRSREXWnByzbjJPkKE/mzpUgRD3hkvHrKVppFckYt0dVqmoq
LbmonSmvOv87WRD8GnlFm74I7jAjt0IRB4zLVsUaBI7xbanEG2dlC8jz48hnKknd
5uxEuxdXHVT1kCOKe817UBXBDcggEyzP2uJDBpnjVBcG5b6dpbxqWh9oYMe6JNPt
5tDqc1A3pibQpR0S4GwdUl/xavKuxHN1u/kPcPjYR/ZoS3UM8RzAPtdTLr72zRCz
CL5YUpFRoTpZcauX4cabqxuCJESA2e/2k61qjrj/aLEFxLILIZIrLSwptByarzRq
OkgtvOsLdLs8gqxVrasZSL//W37KPVuY2um9tXtf5z0jjB5JIDNgREGDYPosl0mS
GPBGGT12R7xltG9eSeBBP2Vc1C60iKn4TCJRLCvYCBSNsS8pzdNm8wWKIh2SmLLr
4kwcZiWx8Zu6N6g61X5aWZ1P1iGmGUHIAR3PpF6jxwFxLWre+cyVU1fQMzjSDZq/
tTqgvlGsnEcEUPHp+C//9Ubi5dsRvBhSN0xZBC21MXwSKtWa3cJRYIBgjbaL9fiJ
MSpFPi4Drs4An/VZuuHyYZI7Q6lSIN2rl7FkMTfZzUkkbPqnqehWVkphj+tsENXs
hJQlDzdo6GbMCMiJnyFDPC07Yq8w/TmUW+i5ZN0IA1j/Ah51HOg1aPy94p+CraB4
VzaxlTQXIeu6Bzs6LmfvF2xvKTFiAxMn8WDBOV2l7Goz/iG1xsmxRhZiaQj2nPzL
r91haO6VTtmzPOjJzEVhPROeU2PW8lQo+468v7McVY3A4+ZJqdkEZeaaxu04Sqk3
/0lnJ28FoTQ1w1rGbi+Zl+minuAmftQ/1tYbgej4gdD4oMuqvu4U6jeuIlmEPbtL
8vjS8mGfg1LkThmjR4akoSVHBqhA/FoPGWMMaHjBr9yAIx5SnNexhsb5NDMKcTWs
WfT9beULE0DgtENxXGD/yTyfRgN7uh8XPTqeXghc/elUJWsZ0iHwjmKd2uHjgdFD
rilZoc82abmB0ll5oPYwzMuREC5/lLeXMYa8H4GpFtvqIKVm03IXcpC6DyrnNsep
OGlZI9KSYSQJb23vIg0Nd+UOFgIJSJNUyZ29RWsn89roPlvSyioQC6/0Gj8WaJBO
Zs0KuhID42Z54UzaW2iUj7kTWMB8E0mt+MPQLjypD2gwRjG14Zie5yTEISNhYDYT
yEs/jbZcHt/i9zDiTVFjvQMonoRepjUo0SjvdDnqOuSWtVcYhfn83dZncTnAoqit
mSX1+t/l6CAzP3iFs4YZ6qHPG3Gt9+FuJCbyuj+pfDKLlF08ocuYW8XhS9zgPbWS
IM2S4+8bKBChsgAFTXG8D0YjzG7xD/pAYHctivZhO8jn4rg8BHEhdUVYlbz5D5is
uyEi7O1tqO/8/NAGLXJ5sIUxy0nFdbtsB1RTCrOFTSPV6mRRj4h0sk6puOyL3m1J
7Mf50F2JrnVdoMIDv19PuEjTo8dxA26rXA38CRj+DhW23aqZShOq7w2nd2lu8zDo
j46XHuGCliflzp1TmZNcMg1zmd+AC7g5yI8QOVJDwKOPR0b3TXAJfbAzTdiJ7Sso
cxOn1wRtN+JsSTDKelEbc3WJue2rs4PD3fHvpvMdfj9jnc4iFJWcJx8eWb05+Pk9
OjoUeElDse4sWMbInIQ1wNlihOgqLwi8PHoZ6dsPjdsX7RAjCYmXk0Z5VuiR6NV+
RqAE3FbHuLq8ozd3rdJ7JayG3uvDoRezHy7rEaF8zAK1vqDGF5xgqT1nLSEEtVzL
gN4ce6XmhBQf2WRluLSEw6wk4kw9NuVsnuyKg2n7OZ96Ngr7Lg2jMAb0nVCsp/hU
kTiyyQ6kGg1WtaPd6ZuJC4LAGGrKopD7NUQE+4nK+GK3L/4udg3+8LKjoOj20uaA
LfRlAp7MIljN1lQtqZnMZh8WPuGCh0VTKSNkRC/hGO9OjadqkYThA0hgWOgpr2tF
WPJiNlvlNJp8g26HkeLQaFF6MpOaoqyYUA6ZMYn4ZUwU7Efx2BIQ2boRvQI6QGgd
YuBmpslabPFCthipZC5wNRnPGl3YxsxQx2XiQOIUoSOIiwvkctH1cPU4d9R/8qgV
ahyudNTyZsEQECjkF8cIUzYYQDMlaye2hPQSgGMPv5YqYbGwTBWglGWRTN5s8mD6
LRsWvfmfMSGFQsl2tJjFs+v36gQ0TqysmZ/HifFXrdgr+kM2FOP2TjnxPjcm/LZH
7ezXH07b6rTeDpgDNevK6kIRjy0YLDlccE1vQIxmVK9FTGnyPKDEFFAYfMzcq07V
oIg35PXCIkC/fkDRbncoTNJqroifLaPEpUDpX52oYhmSKkZsC8+GCfA5kf1T/02V
ovm/NphYrEbnKW6JtE5BJKE2hf5JKYXd4rzMkWZ4gYdUOugV8xY4WN4Z0xu4ir0h
/eY5io1E+6KiPqANU5WHZB5Kdi+X7Zcv/wQRMyyz9FYwEbeGVS+3x6aQ0GIObogG
A5tu7/DJSG9xeVq010sXn+LaqYt1aK8LD3T41m+r1DmhA8lNUfEBI9aKYQ0iCvc0
+OuHj9TBNJXgy+O1F9KI0CsxIw9+ypXGqkuTwMe+q5PgadJ0yW/GXiv9B2kE3EBH
46fuo/sXsz6UZEgMn9y8GPaauamhroTOh6R3IJuiSD2nvxq+tHbeV3V+9l/x11QD
FZy3KQztuRuUABpi4TDEDvmZOaZ1FU6rV42FmeyPIOBlnkHBMX6n19/TKNPsGkKo
jJQcDz+4vilQMolGmKvxK2lwcLYaZXp3iJQR/2JDC29vkCt2vhb7Dh7ObceeqgpR
sVCrvsqKp6Js8Y/v3LR0rgtIFp89oHJUSthIgXioExmGuAR8Ix4PB1MSfqIoXx/F
qSubGy5ynbvHeV4+yC7ws7qf+X9fQfZWa1k7Fboi0GGJd5D6VDKxZq0J2mT8rVRq
uG3TJicw3qGpU7nPyWbkuGtVWOkR18y5nZYtsL+/zlotF7cN1qNyOL0GbU3cXW+G
tx5/lDVwORrUPAY8lXs195tG7K7/m+htFSztXZiIp3y6zMn+1aGGjqO8GPDxE3tt
nmDO3+19VNkVqWdZi+oh7a60PQYC4ureGcVv5+tibDTK2drFKer5a8g10DZkz6Vy
mqDm6z4TAkGK3WLfMlgpjptPF7cRKTHSV1g1LSD/INq18B090kVC5AC3+3pX6ZL5
rArHUnwjb9CRnuWH2iYg69OhL9hZgiV1kuc+VQxe0KDDQ3Bo6+ePhg1osN5v8TL/
VxK2QWEBac5yyKkHlAyzjQmfl+ZRVW0KyD4CCeDz4CKKQLuWFt/6vFlyo1hoEDK3
BcNN72wIYAztBnXYTx9FrGYcklkUbRqrm/DxmSP1+4qHPHmCCTwRbYaDyyNgEI/h
SmsLRroFC7/VQxC+y6HT9mI0Av+5XL5q8gg+/lpXpiG9MCvbylp1yF1/RcPT98VB
SQ3GUyvOPhAixRLUFuRw0R2J55AfditqyCDLmWeZAQ6u3rzMrtmcWcuT+v2p1qrn
cIMtWIl3Iaue/ulKPeHchLekyiy4cn5RIxUnVVM+K/3Hiyk7sPP5lrcJTfeNJf/M
mNOGwjoW4fCCPgRKKqF2+dFsIBpVmAOpO7ugkOaFWR4zrNTFtBUcBgUgDknLMn0S
P8vAaDeI8EOnYa14i+ZV0KWs+31I5bUfOLT/WO/PJaHmgjkdtZEsi2MqsL8M+e+l
1+8ZsRqZtKsPNcSU51eEEAdRa7ZUy2l5caI47MloA0Xn6dkTQ4dbXeXpS4vYe9oe
fZsCefHrctjiN30az3kRLx4n0TgLmMMs/5DC69PE6qkNSaeS1ic6GLBioKFJ82WF
SfUxdFwLvcbSuS18peQ3oAf8dSWLZuK8Kj94e5fh07kn8PRIroJ+VpmXn1DOa42b
pBSYwmCli45MGLOtjqqUodSSCE/tdvDVcUybLHs6tcDXJ/ETq7fS1JbYSuAq5Pbt
fEaR03BgrdsMMzVyqDUwhZK9GBjaJYCDEzN6PwDIAk5+3bQBQ2Rq+b+N+PNPB5hc
poDpZabt0zBNvv6vld+5aPlI9WhQ9wH5wYRtzHVsOJlcqLZgqASBijn2ipdhctw9
M0LvYBN5kiT3geqIyqIIrkw3nHSDGDq7VNd8ZKhnS1ZLn1+8VETPzV/o98hyuyfT
N/vjABdzs/K/hxPF3XC8VjHKZ/I/115wZ6hL3hbIP7pAPqhcyy1QzD7sY37TVMAJ
/OGpJ8lmL+dRwZW7pyzi1Xk06DRVjTGQi0sVgx4HtjDIn66ZgJcP5IH6FL3oPTQ1
0wOZYuVtI9qSxbeHjTK9Th5Kdvkisr8kFBFRDvAfsuWISlZQSeq5AWg12i2jmGuK
r5GwiJal7HkLQLQDrLgp3oEgFf5vp3epj49qg+vvwDpR8v3elYqU8ZbgcA/Yk2xl
R7h9cGZDQ6V+qWho1mdGpF+OgrbKui9kPtG9T/F9DoZMt9wd/WP+m/OBjymGXZrd
n1A59cbAdnxIdcMxgpxM5GQ2lvQzWi4eYyfTJenM4wPT2dEEMqb2tGZMk7EfSNw+
0pKNrHfLimvmmNsDinHG9eMN3L2zcrbtLGpZAltbjMlLxbJk6PsE9h91QwDd+7VG
dIVbbZPmbGxKHUSrcFVqAo2pAcNsPrNxjzOr/yvd8NDJj69rmiKyXYERza2yKDNJ
02+yAud5XbtjSORt9sklqOu7s52Ogur0QTm/XFCnozEk7Vbtdze757sXya8Rr/hc
pZTW+/Y5tfMY8au4WfDtWiDuunkQZ0nUwQsUUpuuIDwjEEtR6s6GuInja1TufHgD
r5u7s3SOipFP8MprPwLb8m97PApl3TBWYXYsyNU4kulU8dy4pxXa52k1/+I+NRcD
6b4FrR3JjPb1riMtdYbfsNpFRe/TtwyWU7hA/qW4x47ov6hXssMoyV9dzxxpuVPt
El5T4m8vf58V7u3nIlMpPM0icTlSuGeobLkU9NEU3xl+Hr1M0G9ou3OAQK0Q+gep
N/Kl1tn3fuoI4v/7cuk4rGewzezTeFstmPigX0w6IelwRhkGoOqBl2hpMdm/KPMs
mJbY0XnuvW38UJseceGpqm9gqlbFkl+186KRYFoWr/h5L9zjZ4Tnd58FHcyD836F
CkmazHCR5Q1w/ET9kzqkR4Hw+VFJhA2/Os1PLdDnBgVJIi/geNYRHnE+BZXK8nq/
T24piKjR0VO9FZS9/ESh//LmcAYYPg4iFUz16ybaBfJ84E49uuPSEPAzWHYbNm2P
ammpTqdGeUNnsewnsWmLRq7pqsrGAEKLHa7kdx9R8q/hSD7AqLlVH5LD4LOvxiL2
AqCEC4qYxAou900jYqoIGtpPNxeXgUFNVH9eqliMbeWwD9YQyVOsFup5CL3v58es
+ccPD/l+hwUQogJd2GbNQnZ33YkGn3vRYRZJ046QGlUZI4rpQjvK2ydFFUmpJrlC
mhJ08vCLKjMeO4Mah8Vonc9zBoE7eki6KWoLgpF/Rt7o7pZeUoah0H43DMER6Frk
Ce8Kyms+xhXbdYqDrmmPHK2NZfVs+Od6qRkHN+U4rVTIGHJI7G9cRyg4sRBySysg
m7jZipSb/7Ou8WzTA2Sl8NGL+6qvnfNSkjozEs6QkkS8603D92jUTJEIVM0GjprU
8dgyxlWVB8RwNRAaG2Z7i1iQr23p+H63Y5FDSk2EGJyUH+le8TcOxcstA2KWGuTQ
7mgCzXUqJT+zTkt2OU3EPw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hd4ifr/awAZ5mHW+cD2i84pQFCdvILqf9jsu9e9Yk73dwXXGAh5EjvGfmUNAK1gc
EEoeyxrOAQ99VwlM1hANDdJy45ezupEHO4RmeJ1fBxljjhXJK/pLvLiVes/PfT/8
3hO0+y4wCvYT9rAWBFt6ToDCWQh/bDmA8lMjTref1NN+Jj2cSFRk8OAVE1Px4h8C
dIWbMv5Tw6Y3MXXhk4QeTHLuRShd1UpXFv/Pceen/WyH2EFgu+GorvaDldAR6G6u
KjfPOYzNx7GM06BoLnUM+7xLKTK7TW0fwc6nwwGeVsAX3tj0lxAM3jDy1h1r0KhY
tcMfWm9cCE1AiFqw+r/JbA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6288 )
`pragma protect data_block
DJKwltJH+tMp9Axa4TFCx28vlDs3QaedT7d1NNNDrACuSu+bYBbsva1FlJEyDreo
3yxEx6G9dg98MMIazS9P9fTtmB3KMZvCFXVBgxkItJ3D4MtFxagkgnIFQuDnFpoQ
tnciF5mvTBML7lLryB7ith3nxGEIereu/vrLBqnlGQ1MGzXsvjHXNwdYJS7HQQ4C
V9ln13ITROy+GYJrKLQL89/mNasrFqYqvOxiBcXb2KKazsyn3YITc80EqfX0axfY
FKba4qawiD+sLV5DB0jXC4Mn/gTyENgxsTMDhQjWxdimwzLp+CqiY3Hz4Z2wixS5
ABw6OafTXrN/SQqcy3warZTpYzDcg0W3jYDzd+Xetv5Um8rj23dd2zApmNbd36ex
niSSR2933S+YpWS00hA2bZDHVdPruJ3nWNeqBKwfCW6k16rr/mfFfCNqhHimg3OU
0hzY8UVGUvSoe61vjmmz1JNJWJxxBb0v7o5sz7cAPew8wIJUJzcVlpidF6aVou5m
+9mFruq5fV/SMEgWcdO/4y8Rd3mBWpehv9e0Fnm67bWrGM0Pcl9FEbtvopxZX5Mp
js/+Za3gwcLPwXqNy5OJ7h9BLH8HO9TyG9M7M1TwjfftB9axeSKZP1Dnr8EWQjjM
4piDTew3YYVsDSUcI4YRlY9wEC45Ar2qDPu0kkEE6sQAQCr0LI0lqx/4qn7XDUe+
AvC+UTHbrcwoTfr3bG6FxaUaavoWn3xoPSaCxmG/lKRidmsFQVJFkkjVNB2LKd3W
2Wll8Tq6n3h5XMtZziORy1yYUFZiLMo9yHW6CQO1VliVI5YLjDvUoapML0LcEyR+
p+28jDi8Iqo/RmVQYYv8ZAEcMpmV2W/Avpq764DT+rzzcWrRQ466sH4VHfLtFTY/
7sTdo9VMI+9yaBuGm/0YtHmbzR0+TTcLUZ/ia3Bhc8zJ13DsPgl/heZL7Ask65pF
vOUyktnvqg93scwlsMc9/yS+5/qQhh4NKVgocdw+Qjph4q3u3piCYtVpojKw9e3D
CqmTFMyXD81xvzStaVx3tppsHcHuO47N77ZAjxIU/EO/H1TPRX2yFxIDjU2PIF/4
kjegKSnjslyi4I5w+VpOBqL1PVCT94B/VpTpQcU5ZoxBroe8QeF1LogxUb8jjMcj
TH7Rvz3bejj9Mm2FyeVCEyf1Rzi8FM3Hx/FDPU1M0nyGcmD7ZbXxozn3jJN7a4xf
7uSgxANBAL+Q4uF3k7E1D2aQK1RSKt3hN5e/xj5St2Oo4w9CJ0x6aVFRNBMZqYbu
s84z15q5hjIxPKroLvsCky+IXTGaVA5DHXdGSRRTnyHBUkcZIQg8aJraHG7Cezp1
BVfcszZIK7/J++V+pulPf76SrdZIoJdO0VV0XBN0n0wafmTCSveHeKlo01+8Bjqi
K+9EjPFNWScywVhitB5Nfb0h/sN5Nf3LWi9MWFQpALH41UubJDnBOBHSb/1qsC5H
OmCyAYoZHn6nVTEuawlL25/PaWDlbeYzTB64n/wSW1Mvuuv+ODO+b3D1Yf5Iqvti
2C8WCGYZBx0N8LpMsFSGRLOIBtdhIelgxMdTvXkmylsIlF9WrMTx7xm+L/TsIsMm
mjf/Fwfy6mGZ7mOhZ2BiKTmgIXgHef/6XA4OvM4B+2RwZaNPLcw+qG8qZ8H9A9PF
TeX3rYkOXT2FtgGlYDA//YXH87adlufgt5EoicalVtpgfirsLJft7A2n4+KnmVu2
394V89q/GpHYcVNTVGtmbTwFRXKLvzVi18A6svcROmahyhrM4vs5Izg25R927FOw
Qrgm6B9t9ybHIjr0LzC2Ny+W/rHhamL8QI345Ed0KCXJV+Nzg5LbnlWDa9sIyyrl
xa8U51w2MZZRE8PdPxTdPYuFqKaq7It+wa2RWl/S6EYpNaAuPh1dd1uyk0VsT+Wf
MNRduR4poFwVp9uSwJE9JfhgLGWFEuBsxZdUY2DrI1zKedEqCR9rSUVtm84xeaVJ
REj+RHdFIGJt4+CtEkzJm+PARRwf3pDP1v8FRfZDav/pASda/8sFeaA6CgzBi7Oi
+9oEy0MUq3R5gcz1WsgO33bSuWrZngMzym1KFYpT7NjRypTmpVyIKlHnRkb1Zhpm
lxpAleoMdwTJk44bG3cduGx16POHIo0dxIB2s9qStbmFoD5o0WK3LUpWQLWBS6+N
pbWmAj+yBCXcSvPiCjenz67ExK094x4AODB0CmQyRENwdNsm0kSD8SaSB9bKOtcK
k+e6BXayBsURHQwFXcVXYKqPdbcZ4PBnPyRkXYweM6pJWtE00M7lpnRz10UAFR62
0rZ4fSyozDdujGfWdVq9z1EerMrIAEOWWWP1A7b+BfcE/TQMN5lfPvxHAGmpAgkH
4SEQGmRe5bGpS/k6tKHe4GQimtbI/ZKAQgBxGn23DEUTjbK35tF1NgHR7VxCSDMZ
PyG4INfJSsJfVix+XD2SZDP6ER13IYpEZGFvIetmKvLDxfxC+5F7XJ0zkCjRca0v
QO2HNalgEIOqDIoAIZnfHrqH6ocCugfSvJm28ZscjByrpEBW3x55fRG6H2Ij+TRt
VHlZ2xmtP295FsxJpgF9yZnY+gO5gAb0ff7u+0afuabFRR448sNX/NpEzyJrMhUv
j1fp0ZIQih3d25bpk09lRuUlEDfi+nZOwb5KmE6h73T1tjF9F3SKdHK67IG0KJRO
clBU3bdRxoLWg78cQkGqfa37ydxGCe8pcju1vdoY+fgbidPwKY31wQuYlbVULVN4
dyAkRMvIIVFqBJfW+cMziwghlm33xDjxK/FYc7zctzeTQsuxV8hhgRn2lTW1mlBC
qGg/WDMZ1db0mlvA4wOb88tOZft/lLdQWdHpmUq7OBZWyLzUqNcxxlX4yX3t1bAQ
A8fZ+ctK+1/lnc5R2iVe3Ozw4hohY3WO5UuzgC6pYfACYmzoHd/nC0csj2KXvI54
MeeWjmHVwqXINU41Bsl3W6gSWLoHTHIm1ErdpI7bQZM+BxeF3lQqnR/776rvGuIX
Mliq6GQME7Rm6i4KIl3uh65zB6YD70DuU3xayfOpt1mjUlnrYendGVYdAK5QkpgD
9OWKs+MG+YD4jvqHw3FWQyzdncZYbzLmKQMGotRf0fh9ZOErzI1kS+mUpPxwO/BA
T6dZoyektzR+By2cJD2/6AyPHbkCQAbY41AtkIDzC1Jm8sraeKAI9rWf8SIuCtb2
hQgO7cfxZnYdnqJiy/hc5c1JgrMTCTVde/Mx8svqfaUiVMAgU86ltBPUOMY9GLmK
Rp9b83vka3paC9KLj0uFfoD74wzJiWCrVlz3GZA+LK30h5qXgOb4FPRO90kZ/D1G
fqgKQE9eThK/NAtv8Y5b/I/iKSB9zKaD4ZvvGSilDZPzZwstGZThv2rTXJQ4ZRNr
EZCiKsSg2aSxKkgEPDqH5sdl/4fgvFbnob/stH6HIKwWKHgd/h23eMKMi3Oldpkt
ROk3QQcUYfuEkv/mZMAm0XVmgurNng8qhhFQhs8TGRV8Vrt9mIJb2JuwLrowFEuB
4K9BCYFbCxiC05DswlD28L78TiuV4g8gkBnc8vCWRCIQDN8Uoc1xWFqrvbWk1/Lx
jifL0w7unAtYhaLbLehOfVtxOUzeS9P1+WZUmX8HqRhE8kDkPDx1Sak5BPuJEuhx
FYAkpGyjO+JyTvwc6QHBYHr/uT21oFu3Sroj00luhVP+fFjkQ0epG4+wg0FBFYMq
C9ChfIGQp6v4Yn8QXq96bPJtIMSiVpG94yBryOeQDMq+gRjgKS09LrJvzbHqrA2Y
ca1xDCEzjnX1iHSEeKi3giUiFLusmrsTPQOCtHroWxEMCD8EX2Mje+aBSPcJeCGa
S0NsJCqnjzfXejY7BMo+mMTCIAzOKu0UzxhzTeW9Cp1bMxDuepVSiuDB2C5hbKaA
eSI1t2SAiTpeQFHr4JYRKoPtr+g54lm2e+AUYbw17xKGl4Kstvqd3Z8XJGvw2j5s
3BRK4rtopGUqcvQK/EdZ85beojlBq6u4H+wZ4YnbJRmHbI6+TrmhLy8979FgBVSt
vM3++kHTRuhAU2ENlgr/GvXvwtDQVQ1gD1g5HmESvd/hWWBISD7IsIaZGg/dTeIh
Rk5umZmgy5aZbh0cSaNpHwVyXaq4PpD0vYSEsGyY7MN4putKf7kExMJM97cNHJCN
ReNIgZnEj14G9d0o8c8f3HEkDXE7MNlAuQ9Oes2xS+bfm9rclF8e/9EnNyOjFGju
RiRXJrLP1d3jHZxwYnxhnHG+XepeGEySxQqGQhrC4rPKutxgnQT5HUrgOibMPjCH
/PGoSoLJ+mGxxS4JJiRYnPyT28RI0KxArw1vpWjFomzDbOj5lisaB4W5b5FGTcuA
BuUCcDtQXa84FlsnF84dLaZ98JEUpDxHir9cwZTBRFRawSzCLnNg6Ojy+gk/u2fC
w+9nx6KI+s5GvRQ5DOgaZCcwYIOxyJGYpcXoAxtLf5DtvR4vrywGmLWnAvX1unGY
uv/+iyWLuy/nNfBAYfs4iAhYcJb748/s6BTOHL4x3TmN12aztt/FMNsjYKegYj7y
52dIHbmDcbq8Ck67uAgHMsAO3LexviQpRWjEsYBgv3DZfVJg6ALwP+QXNTAUgZyr
VGNww2hcpNWbsS8ea5rZgdmumpPPUTCKkLbT/MmiNGc8UzBVXPqn08PKJIFIS80v
z9Khcsl6u0H/y4cvTalhqHKCVkiOMhQDSjqifCLOa8tSJH19kv5yU4nkLu/PxP3K
+vdqbH2H2nM6o7BWaQGoV9VFhDKeLL85LB+NOROXw3Qn8xMKN/ttCAk/wWsenZfe
NbXa0y3sH91+zrX9/VB+0YVmjrIAO9XcyI6yqTMdUcmgcfqGSRH4sdM3VePeHVlj
Fm4EeK5xZzsuxAIR9SmV44ZXdgLlfGzONmZkvLl+A450FYjsfpVPYXrLlFnDa8CD
4sMsb1ThmpN+yG+QneRwjwrTO0EWJp5RdU1gfiRi+I6PU4WEMmYU2jB9v+WLH3wy
sfh8kmndXpDPOG6AUM4x3lkxFwH/LQp+Q+QHGorCbKYySNWDWD86+GpvamTVHDID
/JzuzGo/SJA+bCAU2Mcvr2+F+92cTpI5zQ7xagcZPgB48RCnN/tu3VteTSKYKKRg
2RBdvm0ySFi+Axbfzzr/e7KxpGZaGtJXEU0MKDGnJFXyybCpGQo7HkxsDtmOLb94
RdbOlKoC/bicM6ygOyKqtQoRNCSP06UwxITMDGobxDL71b/fv2v3/xmucYUDXJ3a
RXv4wtY7lsUGgE00MEz+E2IGkNOLzgUQr31BZcAMC5YebK7kGZ4r3LeW6UNngGJC
IhzTIDfKO9SATQdneFQVRPES6dyz4h6Cy0XH5wq8+MJdxFRBrJyILZ0n0+b5nsh9
hQtGzplMyNFGgfxmJGeKxjI1WLEWym4c2JYgIDQ8oRHzKt8DZuzA8nbn3J0mFYgN
dvvIWS9ipQk6t4rwvznPR+EOQVApAsIKodoL3upAVmKXg7UQ43nQ97Zy5hiCunPR
i45zs0B5V5V4NRPZVVPdonFpmsZLlOHiCbnRUxHHP1LsJdMSlZGaAi5dUKuC/1Cn
cbXz4gYFTe+yd4isUDw74BrcKo4YgDnTn0b8JBLjbZrQa+bn02mPG5M+UP7BdfJG
1rLnbuHaZmAlJ/2GoO0GXK35Egqn8sfbgKE7ai02zKMpN6JKdvbWBr4fRbmTnF1B
59ss27G2GNE+pJZcS/d/3bQz6Mi/IwCrZllVSrbLjKIPMNAS/j9fi5dv8L//66Zj
DJJY4BsaN90Nc5+d50hxWSBdgTQqifuWWMJ1M1s3zabsMB8ValEXWf45LRMeyZIS
HIPMwc4O6uT+UJ4kXxeMe5O6RlqqVgTBO0uGs42hDQGAcXWXdHizFEwdzSCrKDV8
zsXdb8s0CoSBZECfc1MI+qhaZtFwTI3XrWmhnooEeP2Q3Q+wt/C6NrGSQf2UOSFH
tpWlz+7kpyDL+bBbijGLt67AZ1MSe+aWnnhdICBUvL1htCKJY1kLs86dVOHvSi9H
I6imXG2pJlcnvA13MfCFqXzGr8WFytf0tgXizdzXzK3qoYk8CCC9Y6YLtePwTOwa
Cu1sDMpHumFVgSjgTfsKxEgYd2oa7stVICqOqxbYdV0xQYDzrwFEMBAp8+Iw9+uj
d7PDr5ioLO/jBrf93iqwS5f8wpWVSEvLq1+HkIQX814KusYisOiOjk7nOpnZAGLd
sfAwlm/gW/oGOXDafpex8qTlMrN+/lt8yBgxHCmzeQETWYi80lKSHx4a9a7KxL18
qz8YiVzE4Yi2JoC4ka7PCDThYQdlTKxfrWqJNs1ITtoZo0JEokAZSNJ9cAwyyDz1
yHk4MOhKrr7SInImMHn7fl4E4twnx4/MacZxzL4l4R/SP92IObLN713VIXXcwA+Z
vX7ksiU1BRASIKgLtDbKaJEYAfjtNf6CzEkCKj3TJjDQ9bjWHw/YeH9f0b/aFiEx
b9D26cEmrFBw+FcImOXULmoCDmKEYJIBICHrBgYcO6quzdiI4ZZNK/D9OHDoxyPP
1x4I6ZUOmKRGEWDzenuPQRFP1mWQbeoIhiKSGTo58Ir1QtSxlDp578FSGNoC4LQt
7joHxZPGDi1tYlyru6F7Lj5Az9k8+poihxXfPz//hjmzVoOyNtsGZTl6jjZckLGt
bAyp0sR/PSorbVpls6U9c+jDQ0RL699u9xRPyQRWN41lLbG+LRru3HxS0uIvCrjQ
sq8EIIJc3OFhdLdzqnI/99aqhF8IpoxdhAF9tPCrUlHcTxK8Zc57qOS54bzUQIph
YvJEAhvMKouL5leLt9eRNSN1TZFP19h8YHE3cnbM8616EdwX93kq30Y3fFeNdG0j
iuUptXfDRGtvNNjairSnHq2HoxfM26jq2nvc814/ekE2oX0zZgFoU99/HOCPry5G
fVILuYxzen7wiYcUnmShmuTH4ik9QkQv3zAKtLn+vkEOK1o+BlnTFZcPZvOPuBlb
mz6o9NhkfaUbdfBI9BmdIuYhTp3ZcS/5Cl+scQ4LDTUxgjTNnnxTyDKIuDSfmPDC
LuKjowj7EeT5ZtZimzKnERJGolziVHvlzh5M2skGMnuTKNY7SYznq8XGzMKE6pQK
+GYq4zohDdH7lFO89lmR1fQgz1oOyNjN5NwTjTh++ptFjuWLa8AtwEX373mqJaRT
4R3l0ofgyTrpcHmdafG4fJSXNKHhXJxHpvuACG50ys7nPLbeimCmg2QqzCTxNEzb
GRiH5FVb2l7X5/qu4rv4k8fypNLvl61TvUZGNzgOjWRcSa9g4zi0sbo8FALuP86y
alRa6pBTcuTlIEvQn6+Mz4VwjcvoBDrb9eM7Kxxx6PvObUE63dTE2UeFr0aK0f85
iI3PVTefau+Tk8n6iEFn9e/G3vPSz7lMRmvkDGVRuEVvPVgs8m111HdBPDt0zLDB
rh3WPtVBvFkVCJsvEnaot1skM+1vF7R8SpowARXTcfBrYbV61bEhjalCCncnvvUZ
NhOIK0/3ztDi4GbmWvOzHC9kl5lJ1kHybyJCtrP0LIOz70wfe/4xLNM4lSFRN/Xf
nZtH1QuaXzw0QG9BUgSSWamTlRPncan+BaX4ke1+H0qJ5RDyaP83mlo4aRZlcI6a
5j2tDXHeINvhKKWpdngLPQs5ytUZz4G0/IiY4r/WncXy3qBnrdrMLu5jTM79gMHR
uD+RUPCZKkQLQulvrWcP7A5OAxXm+46meDx+MZYnpm3k0ITvXeFsv8mcCwiksckZ
rDK9HaNgh+iL4/oIClJTp29AyYYmr+YgIIQwlt/LcGi3LVoAsRUgja/a4tdWaVQ/
nKxpGHJNBoQ51Qc1jlcsk9s5ctn9tTc95Pfl2K3b90VzTRRnu6vn6yQ4lYBM9PRN
uSFFXjWxmZGQdWadjZx/S1ZaJAbZCsknx1r2GDOJWZLQUywdOO9/Tav2x57SErVO
MsKrYF/Yw7OL/dY2I5cAT4vgqNOyKb4WP/RKwYj07ofz22m187chSs8/BrCx8xVq
Ko6nToJ8lTN3cpnNYmvLgLrkTp4965AnRoRow6GPyn6anDptJw+jm+Nj1rqAXT+e
PrILQFU4OFZIAuV8T8NBOhT3IrA26OribGfo8H96pGiIDqPjCVwv2x0jKpyzSwp4
Xsuky//CM0eqqLUCvW87FZezlzszqSVUlucT+g0BCYG2xqR17zmfuHqTtkYFEOH9
O5U2INuF/fVSEudoFyv+Bk3PfiM3OgwHQ4D4XB4Ahg+2wOHA4kC8fpOTgvtjQ2Ds
KMay13hxxtOBW7BPSKsiKoS1vZ3nYRV7cOdFAF0oxCQdvPjUg34AKn5GrdZLmf17
rtGXKdpSFXXXRoaQkJMEox/dEIh/GTTZpScT5RDEpIS7mvQ6pGrraWL/DZPPertK
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lvIdgEJ9RYyLvf60PQ0XoLdaM8sedLvfL8YLK07HMtMwvCsQwKHrsxi6aOz4YIky
VpAxQcFd4a8DClh3fS4UqgKRW6+HRDJ3keaOmNzfE0JmPjDEm+ABq5JBhxXnsA0X
cAcNwvjlCbOXfQAdWfLbALBDzyPGqVAamYRgMixt8euL32BLhRwrBRceCFtPFjt1
pn9kS+gsy8UCmk3LfSSdM9KkYSZz453rGJbcP2VldFOwzYOMmu+Z7dMcyEF79IsD
RckNQKkZ7WSDMTn5Xiu0rCq/znKpKJhiBHpToR7aMIMENVe7AdNu5Hm2+VgQ9jGM
YV+sHRr7HQ++e0GtVAQS+w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2496 )
`pragma protect data_block
Q0tEiQkUCOvX7MWLb9r3vo6WPUZEaDkavFjcokz5O+fuTPp3vXJCbVN27d4MiBVZ
aRHtPNPc1AiaPkMiC1WWxnY9hUnqyymAYMoZd/BpdkXKuTFnP4NUqbiNhJmuUhMa
f+YFkOqyam0hDhS7Zp6KSUgP7wXcP/ssAmGFFeBTbjfi9/xtLN1RXiTo+VRTCxTZ
4ojU+b5zwo5dr2w3r/oEXIpppHkC/YHmckNTdTL4MSzcbICeI0QWtPIEHU5xpTUy
FfVh37UeDLqPu7T+0Sd3/thgnm5Zvlh16ASlQMbnMvsYg/fwBmMD4wuGZIzjLCS/
pY/zEag4omTfUpNr43auxT0NVQ2IQQ7viCwfMzwIHU9yUEVEQ1Mrl177/BDCkNZZ
kbYaESp9Hg853pI3ZLHeiocGcZJh/wztzE3kbNMHBwt7EFRFqwJrUYTKZUAUrUE/
/yZmdEA19Du2HDpOn2zSnRRJmbP54Y40gx1BaoujNqgChirHpjhXdKXzIhWQSqlV
5VjNjyTVfxOcjg7Z/DqszrS1yJ6rDoQXJ+OzrX+YsYHjF8xrYe3DnPt963ae01jW
rrqlNDJQDRj7M86XMnnAq2kaxHJ0DJP4VfcooLkzHAbQbiyxCppswRaqrEfxUYrj
qMT3Uy+4Tgh6CcgQmuAwddHzpg1U16Q0hZv2TUo8cEIEhZdCaUAD6ITF31aF8XEA
Jcz1cQVln/NfF7GBlssb7CjSGXCWu0j1ot/5Qfz079vjVylkWGMdAkoVme6/7dH/
JhK14DgVCa8htosQf2ZD7RWuSXRBy1qKP8+pzrUxM9mQfdMyH6iaeK1v+eD6A5WD
/526UOuHdTOjy+XuoQsBUiTq96/Yduov5rCJn3wPAi3GEcPtQB6AAD3kfPv1cV7j
TQglOiZ2j001sjIEvgzcsNmFEDskWF161zG9R2qihkeRcEr/aBnOZ39nII3Ya7vd
I+PioIvyA6Fvi3nZ7hVh1yEJgse0t5tJ6rUqkxsKKb0Pp0dk7sPJ7A/pHiNY4AX1
S9O0p8r6JozyzZAq+QUfAHuO0re68fq3OYXttGqeVgDC7aTglwMQOxo2Q2LZQoNy
Yw5XgkSlSeMcWB9NNj7YT7wUxlwH3TZYG6il4reLIHTcVoAv2LNqOG2gs2EBKsHL
rkJGgX2HnF79sfp8zJAat4oM1VB2Yg9OD4UvmRfhXiFHGSypNMB9+bagQlXPcibM
v8+NJkogIbHDFFtcVntqmySTwQS/VNey/RCCucr8RmC5LtJafCishDqN2UmdVaRM
0EiTOQSN+saPLQ79FxKywodWwtcKyMpBkVlpVBEgL2VSu4nm778sBOtCTkIlBoti
xH4dCfMOZcmiuCZ62cNDVVQMiMnhFjotMr7D+d+H6REcgo49xeDXAYJWBU105aK5
hiUdZrWpS8XZVY2/8JMyb3cmeu8p/DpqM0uBodFbTPbCT7CLC01Yyy967zO7P2sU
HH/ZIx7C7j+rjCXkSmC/Jtblc87eIvE4FisIS2UJ9Nlr/h6CVf/6ZuIknPiekmuR
x7RZskkjrnGFl+7vLvUP2J3AEPkcv0D2ZLVregTMN7Pydg7WeSMNYF02buVFAPxK
sgIw2stCVoqxO/S/18aKOZusxMq/fmXCIjrLtBU5NwvG++648MRcBKdq8Bb5INfA
rRSxmN82MwKf3OdyscxEzBxIOb+oKDUBHDQ+W8OpUTeqIvmF+U+CmtdXBn66sOPW
f234x/+mvwRYrau+T8/2cXJ8iatHtTn/PT33VLamDcyW0hoNHKQbZn9PztPSuY9C
pS8lSYqYbW/6WO9WosbDwHRruyCF+H0wW97ZaytIJjRk18DbYoAuFNlEVQCXiUQ9
sHHvo0oiByfAZlccVLWrYOHYqNVOynYnuHZCoKoYgDQ7xS/PrMs2P+Nvkh6p80M3
2Ug9vZpSvv5HwegbTy4RzB7riannV8pt/JDJG+EVpZlhQ9IOkIJ9xPqKlSGbJtMn
vS02Xyi9WMMle6V+MALJfyj6Wo/xKiCWJKav/Gwy+wLBtmiIvI6bf0SA/Y0cUwwP
9Ol1ToqhYHtJWX7mFXun9es3HyQhsKbgzmcuTVok/IYJzsq8LULEEqpQJFTHUlS0
Wm0E5oQtSe1/xE/M9/Ys+bLwDu6y+q1jOeahXLCskrV5hCfpthXM/2e7ursMCxU/
2L2wpzqnKkVNkeqJD1CMbNSOiCwmVjLZCFLYYJewhNUtNKQKBDqfjvgGykD20BGL
EyN7Rxgt6sUOQ5no/U1T19jt7ULNdPyYC0eI8g3iIp4RYCauAnlMjZypD4SwkDFa
41OsdHnz4TINQgyHBAfGFofdULUMJqqy0H1hvxO29wMTDe4FmTRIa0ssSUWNpt3p
NtQnvabYUhjKoLQhT4d1cyLasPHo1pnz9vqgiFD/cTtAAz+ihTtbuvoDqHoVUS6f
5ACH7ytrfKoz+tB7BBurlmJAwgO+cGd2tLvUaM2P9TTqc6yRP/0Yd+4Ns/+LvSa4
cN2q7w+5m8DHITP14Fq75+V4oAt5W9izze3izqnlS0whjsRpdVCDRA/e1kt5X4EE
Tu/lWw2r3cI2CFZKtqZLPXRz3H+fPlvrHGLiifda8NFOTcMhi/WpLpOTzYRN8Zxx
P5GfVqolGa2AZzCB3il+V5Kh5IIg+MQdmprMabeFPbf3YzvR29tHuTpfwRxk4zY7
wdHqwmZVOSRd+izMCgHsIh6K6iSyEUrN2DnotzJMnN8iWGVfsv8cpS7qO9P+Hvz8
Fk3vEzfTSLB9ot5jnCtSpUiUzgzj6nmMbQfFRH1uiWocoFwecawPHywVV2xJP9uY
pb90+ElT+DMIJXsxrhruamBeEYhq050YU0phecWRQgTYxwD630PHjWiQpbKt+7nh
k7Ln6X3Ufz40394WFUy3RAXeqjN6BEGpC0npUP44K5gFwiWmNcuhi0RyFKY7KLr/
J9votEvDooH2NTYuTrOqzo4QKYF0FlBCzSjWFJ/fOmuZgRbKuhLt2H8NiAyH/czk
pszSVgjA7Ug+6Cq6o+xS4GKT6dVs6zOTs3q9d+M59Z7J5WX0wyb22eu0rN72PMT7
NDysjtaQA2p1POaHJRh8QbvUWGo2ZcEIRGT1DDurp8ipt77tSmlf4aYmO1p78L+f
vNZGH4sHougjDwPOBGAWwQi03YTUOrtRo299O7rU7M5vOFyoO3uj9iSxXMudOCLc
DTXM1V1O8bVXSSNucVC21f4EiFGYeAjK6aie10gi6omw2aosZhMzQm9ltYJqz3ZB
ZOSKR35WDXRi7n+L1FVBmcC4jXKW97lq/iyy3c0TbF5cpJEogxt+U/b7/FxYkM5w
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
h6Ajg4j8ZXkewJbEvrBkUl4Zx34GgcW/2VfU7dh7i6PV/zfDl0Lkfgb5A2CACLLD
1U+Y9b8VtIYDbv+N9MS3KrwTVnwKwLEqYB/WPALjVaUT+wb4H2ZRwxoVym/XfAgX
f/IXJe3NdlSO3DoFMOaSMySLotmmghzTVp+QXfA054Ive84ZqX9GH/opwP6TPLLZ
oFNx8+LfU7TVd6pvfZaoLZDTP+uyhfJHVzN/vMOTbQukoroeWRrK/cairGudfDzX
ooFYqQVQlRdlM8S33B/8IU5bkWzDNZZr+w+vpgx7+VBMGyKkGZRu5DeQeB7gSlsg
9WMf4bB8HrSp8rfNJlwZ1Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 54720 )
`pragma protect data_block
DQelDD8FptNO15UhN+eeShjOohuW2u22pEhCGoXKrhaBvSF4ZecdnqC9q/q6Ih4m
g9vOj3vmzDN8ur7VyXJSUMeJhI3cElu0O9M0RUwRJ/iUVhEX5fdf3fKD7mk2v8P7
TPSzoagkKeqqjJ4twLuWFqS1uRSiCSGoeatglfiWHs0MteUyy5lve3vHEuEtmnC/
h5KDKY2/4gpf0CYr6SJ2NF5fn43JWW9dzzKbWn0fDEQNzeu1WjkDqELIqVqRL3fq
jEzjNbfuarMFuhTkT8oIY1F2E3RCO16IoeDLifS5xyh8c6VlMG+vD9qe04voYjQ/
ZnyJ0pgd+yNB+WizVrvkn0RouWgXG+B7VcgvGnWEPByIZf8vK4RE1MMq7vJ2cXNL
hlUXhM/6nxKAPBPXetPDIoP3EAntZhHjTrZzrIMCa+yFaXbFGqiC3/qJjDQVYnH7
kd3lttuTz3ZzzW3BdwfUdtSYNRHx7s+uxnWpFvWEtySSl/fCY+zIhKpjYa6XAORE
brEJO+jsPaHo1vHen7JfBc5VcagTcbatCHiWgtS015LhXnLjkDAn/Lt5tPgm0U1W
KOaGgKb2bsSFy2RN0kXpzmatrMjdhZcECeZCCCB5oBorC6MFlmvjqjhhXHQrICCO
Hh4NcPyCNyuq6i6KNbWGqnm3//ZRE9aXeuAEvM4qdDi9cYBZJXoWLz+/VBvPF3SC
+FgZz9A8cOtkMLS6QNMFg9n6B7PHIl4YJyneDQkylM6Gs7zqHaMFVrGiYCW+M0mL
cQARM0PIUI2Bc40MaPeG0aBBC1/nxtYo9o8u6Z2sCVRXKTPt89wWZQWQBhxG68h+
8yYvr3A6Q++h5gVzNZ+juO7y7jimg4tA2Ck94XHOeW8wp/KToPnIH/ySQHa1nw26
lgOp8qAVUFCOOzCqlH9B1+eJ9l3v+e5IHUJbCiuM4doTUWKWYJQbaIiyv0rB9gpn
UsVBuss7c6rJCZmlgckLGAVP0yl/GGzkP2Te/9k51FEqGBu804DSrtT6WivjgxeC
eVvGSdUx8kqvApMaEXslOXkvvhblU8JxI/u5EYmR5+QG0SJw8prLXTQAqAISgWfy
dmRr7Wa1frWKzmlO7wK0O5beHr6t+1pXtJviTpxF7vkpCzgyogUJHOjqkUJ05Xy+
P0fHr+cdy/c5uCfw8P7QM+0G0KIy03mUAfU2fbMPAd8MKUSiNJASabmiWBPXyg1K
QPqQZ7tZrvocpTNNPtzi7ULsladRoEN7tVfvf2OO7RSqbppNnQ8wc2acQSLgFEgu
KMapkxkyDVJ51leIX2qqcnM8DzLyGqw3jBUxEdzXicc+3TRuT3nEto2kMwsGKCKc
lKp56GOyrZYBmQDtIYkKDGt3cmQ0yE25Z0DTkMbXWeOF/t3AUrTCJKm5zqEDoWP6
pEOFDjxv9/Qnb39vvW1e/nj6D4ICuv2gbFYMfjULqGXu4nAC4m7Yynv7I2cJj7vz
h7PiO9IejC9p01DduYYQ3DpV1FWKN8FJoem+l6NaBs6XLw27hbEO+7IgDLm0b0+E
8JReQakf0ql28OxcLJwTzlwH8FEHIXrzrfzFdU62BmrA9NThBrWUy2LaTR+wF+SY
OK8Ipa38KrX0saeSLP4QHSBkmdu/xpE1KYJtB/XSeLTlNTxL+Y/cPjH0uA3tVAF1
EXhrt6UXkHc7nxT+fvzzJ1/3/v8A/cSt74QRtVfRELeHK4WGwvSKPblK+f65DXDg
TztuSnpQOa0fKcfsQ8sIde5xnsgWbt/LNywjs3PglSaTi0kT5Lf+76lEDJ/R9oiz
xfqAlOQS5F6Fgpd04KPxM5Nk9cj0J4kCIcUh94k6lsdzBg9nn0QU8pi8Fk0EKhxp
vdbQYIhtQpEgaBnRvNN+okjuNlqcIGzcBBD4ueZXzD9BigcEh3ERESRA/koc2QN5
vYGWLWymuLSbvkpeR/9irtLvi7D8iTBymWa+dhHlexfOy7+4SUtQs4h3Thwf4FwJ
Kn4INzhnQb6r7h8oJHKkP7msl6U5HU0VDzKy+mm38JrV+PBPvgWVO7UkIAJI5lLT
nl8+J/SaGmlIGhuHYASllG0lSZbEJVaiTTj5g4jyE6JHsf7QramX4fkYLlsgzRf5
3j0gudVdwKxpXp88t3pJ2Vx6lO+XdJD1j9QfPpCpK+rnuHu1CmEoyzukPoxXy2L/
s25qA7GoBgwf7yuxt3MfIGxaBqu3O6eclRW0XiHGaZYb4KNKNG54DX0ouMhV21PX
rgf10K+BOrIKqyG/1No+UjNguQgWh4yYDJsdf525PgRi60IU6b8DudrkqZQltgnE
NCBvTY+gX769emUCMM6rzGDei2dVO5JeP5E4xhFqHDUJLimQuwg+/bxCJTW/3g7K
JX1ehcb6E1ruRDpj476cRBBwkOOVA6XrpepAMgq+AHVLk/NR0x2c1xKfWVvsfsLP
oJa5OhUmCYOFhb9rbsXLfQNlyLnOT0pz9XV2WNMu4gweibhAw8jgEjNcJHwTWOTY
9INEcMJT7Cmfx6WhsIzsiFwVognHTJTmbR1ENyWd61cciDYQkWYln1eM8mycYTo5
pUrQZ2W3yFxxSU4T8xviSRuVggmGTtO2NsxmAFzv97YN+qAXpVmdxI/TjfVmjfzs
obZR979miqBsCcT/LPpuDEppkA+FCYpzITimnU5t1zcyZxtUYf7HcQM2MiTW7RE3
qUQmdasHZiazP1sUkjSC3FtA/+QsMffFd8AcWZZVentXpS2kda3h0XULESSz0i2v
SMMP/v0UnSylvsgl9eFEn+fHWBqPVoIlW2sy05vwXxrHPiUNb6TjBJqXqHSqbOAH
8LICz5oekCpLed7n8380FYoXC1fZw9/E8m/zusGnNZRWzd9Hm3SjhRQsihxz1BfA
FQoVc55TVDLr42g3Pfg2/6Ihs5TV+mkK3YTterNVoqfe4/4IFewwWjbZ/CZH2IPW
xI6GIXTYDhaOKznsYTCx1qwsxtZzuEzAkkvHwS2Qw7g2BjBPrtn+FePqf/4x9UUo
aHynu+K3r9h1y9IYnZkSVxlQyGyHsV4BvEYO3MFAZCZFNWRGsM3vwAHKW8vR5MQt
7xOzI09OId0Q6o4UrrIajPeC8Go1RrcTIglNNZAgOeR8mzqr+lV2ZYlo4O9t3W5r
djVPE8pZ1BnksP5c67tNXNyULNLugUH88QWwOW8GvT6I+kgWIcaDDfWye+97hTia
1QQJZxxI4+aahPEDxfyAavM98BCbz4QnOHYvnRIIoCCVA2259UQhhHym6zYbPyW+
iYxNBxABRPWTFZdp8p93jQBI+hl2LXKWjYu7efk95HP1c1tGEXE/bAeUAm3Pjryq
2Bvpo12bdrgobAzU92Z7MV8l35tcNF78/sCDxEfFTQKC/WX3WI3zz04VN/Qkzpi3
jsyLAqBJjIGhOkFHmGdtnRS8xuBrtz5yWy0/2NLFvjIeoZWtIg8MU6r+4w5ptOtm
JjujWfusHHvipHppvYSo7OTOTBpHHfXCwimp8/MbD+xGkLv0tZ1tW0ygVNJpwwz4
rP0AuBy1jpA/9KzPMNWMRn/rKiSvBc1hAeyjO1KsVciioHnMpOp60q7IdrQN/998
oUaIGD+h4Jwo2V5WqZpvo+Me7Sy5I8ZznGou4o4gHtzvk/qkoLRhGB3MVRhnrpgu
iVhX6hG69f643BYi61mbKRpvNdwFLKhhU+UYQN1mDvK40RFaHs/ILEZqu/fT2mC0
f6upwfF5+MgWrYsIZCWOa5r8fQZ1HrYVIirdrsGs6eUJF51WjCewZZgwZTR601o8
OX0DTjvxm/gES+0u5NKiky52pEvakJvJ/NC/JR1iMw6DGNNesynW+1N2aL53HDYY
MitBJOByxdxw9vOnBza06O/k7VqzHMegcYq+rroWlMXqYSfu3Qm3DDohzxGO4vA1
ZG2k9jO+OrTxaB8Vf+SVFojo7aI+UZT+fTIM8bjZa7jvZoeclEQz7uHsP7LgvgWb
jBPSf9myrDGSyx5EkxeyVTRkHNpEMtLCvS4dEkI1Fq2v/3+tiDd0aXOenUxYVCPS
9A2X34WRtSjCkTGJFH7AjfwYFT1RaVaJQXxJxB/oMqwOBpYOvV2qKpY9n+xx5VzR
3nSSZwypCimPbEK0ve/nvvqhOaCGSN3zufh+c7p3TOCfsyYvLTDi2Vu6iylgcAoK
8vH0xyrYyIaJNLV9bP11G/YmaEL/R3jwsbDQK8nS9W/bCHK+53484P2h1XSMUvPL
LmGlGZjIKGjZHH0x8SwXYq7C0H7maIYm0/4i+Hi0FlJgTHmrLbX/NbhyR5RC7Ihp
tirxGaxZnj9uCK9XJdrDS7EvNE0Ea8fY+t9jHuJn5EU8m1iOsa8QUGrpIr/f7tTP
HdXWAQg875F1mbv6eVTJhtoeoR+GZcPzQVx0XKe+6/qKeuc4X3l+kEseOaetV4aU
wrxUkqLzLtEwqH2BoX/Etg12hAikvfIS7G6XkpK2B5PcfF7opJ6nZ3+ocA2W6lLL
PjfrLSZ4sD2ooNrWUkxntnGMpe8YYjNqC4Mr+OslVA/87PaNi85DxvQZ43A+Od04
ZLI4C24m1tvhHQ+M3H3PGSxq6mN6ld6l9VBopPfP8L1u5iI+Pli1xTnlZZ8UmDkB
PtIfIjw7Ar4QWbmcmxjXm9pmRecAoJBDDgYh8il2O8QmhakdoyOBxsmiwwvWVUIR
QMi8f4jBeQE6risw01rKzeMjJg9uZo01uABzWMWKAC0OMtW5Ft0H4ed3hNiPsa6p
RtTtIGnLAVc0rkmst0J/HiUM/y36972Itd/d1GGrQZLcr5OrHvrqccVUtZsIh4L5
racb+o2IEX0aZ58UgwJJPPmibGSGIdqRa6N5ZrXDiBT4ERuU+p6jCYF5wcslNTZz
UsglXq07ZNGp8AEI1uaEjZfYw8frIK2DaMeSiIwafBtPaCu57gJa40fR3HdWWQUG
swVkQUIo7fgtcIS6BB+i3PlMyApn66lP6WR5NUbxOe3sFD4s8vaXEdDNzlCPXgxb
MD3Ywz5CjyMss4PcOUHCIiTxjun5ou3HMElgU7l4x3bjsp3OgZM0pX7W42e8H0gr
MLs12YVDnSHzMZMnSS0TQQWITEvVIH5Zql+9+X5shbJQ/ulSJ3+31yBBszNr9OqT
zQh/pdt8Y326OHoZk5LMxOU2SL67dsVaJNeaizeRTC0UYxen8iuYMcARCeF7o7In
YEk2k0nylkeIUmg7+Ud5vzihlijyBhKICf9TDWbLc3gM/8isXFWtkPF4G06VAM2P
OByhJWu3GSZIYmonehBgq0VVnJoZMx4Uh4czqUtQ1zctwNHCBhgFaTju8aYO/jsq
CiH/pge9DLRxFwPPThyyM+2KwBzIBFxFmw0ccVZdnvLHnoSKE1V3/vizJWFSrkJX
gelpKC/fmsW6qtWdWPdM2z1JDd0fIlrk4gy0dpRKmS2m5LnLWRYxHV3iaNaPn50P
lJ5T9oifG5N32F9sbM36Qr9ueYhJySmNsFVzYDdEBDS7AnukpTjYTAZK6ziVhjs/
n48lMCdO4KhETIPEIW+UV4gMs61yqCaWGrMuGdYy+NZT0l65Tg624tQhzyhWna2x
GY5HplmVWksuCqACkyKTz8Z8eLP7yoiB11pdhgeVAXr+r8r+fsZrSPeQGXcdc0fV
kda8s//BsQr3Uz9roP1lnCjWr0jzk5TG6dOOivXXfAKgGpAi6C7SjZcggGVwKmhJ
BSvI44z8ZupLRKmZGxY2bV9IE+6/hBIhhm3dPtb7AUY0dwOsuPhK5S9FFzCRRyeR
t9VUkvTtnkOJYbCNKwHqPNRoHlUyKN4YH4yxgWId0KhafrEL/oBxA/ZsvEwsS4P3
5rUokeSNUA0HANq8vjjf5TMggawZcIXX/N8/yr1J7lSwxqVh+Ix2+gRtr6infR5N
pSVZ+JOtuqr+tP5MpX2iB4cBdXM2GyXILIJESX6523xdJAJvkemgb2lIJsyiXONB
5NF2MzzoCj3mx0Q4VJ9PJYMzOSHfsucWq4q6CaCqRm7XDsT0pw8ssG0icBFvUDVj
2MDIyp/LCqQ3uNi78yIWi3jj6sRTfjQ1wZlqTLyQDhGxowEd7lCpr4kvinVyWzKo
A0PxnP4/jruVASIfoSFHp8LNjVQtI8yyqYQGrc7UY+bcB3sxmKWbQnv8G3HVPhmR
vUw//mJwNNFj+rphcvR02RV2CB56Dw0mB2OtQkmaPFjYTWXzAJaCHkmXlOVQMPrR
iZw/wfo7Y+XP7Uo2fzcDWg5Dw+nnLiDJ7oL7NHXUW6Q2MdgItt6ZJEHeGY3qoY+Z
GvNsaC0L8S75STA6uGokFJMogfH4MVxJzZyTy51tiFhE/cTKvSJ3miLzn6XUH28y
941h+g0ot6drqw+A7Fb1GBZgUJO6KeJxa0i6dFCiqR7WeaVlR+k44VNQ34O26w+H
qQpU6GpeUKgGha8MtLxUcA+xUo3lrYvxVlN8RqDuiwSf7ox/F/Mp6rzWGO0SiXsU
4veIfGNfziBSLml1cLgPX+WHkmtJRPLzT8lOe+OB60srAgxIFpMKLsqIMz9jt6Au
EXy/V8HMoR09JKU3hfNZHiLEkbAmq3wx3mbH8UWupZCZP7QxZFPnefhCQrhwecQk
k49FIIrN/UOwQrpBUajC2Bpcd5A1H+uAq3FCOlqauvxQOzd3WpGbbse0/FEhNrPB
I8oaKqIiXdDBl3NzHyZKJv+GiAMhgQGe/Jyea3dCvt4ASphZs5HZzEVVbglqkJxe
htrn4aapFlAX+eoJMZcHSw5Y3zKIkDDKYSpZ7x8XVPY3paErAzQtZYRWJdCBLRd9
Rg/V7og5wNpN6dTUKNvsjNRyB3UejJfwifB3TFYHTLjMDRvazRTcbUNa3gs4zifQ
mo61+bSjeFp0pqr8q5ibrUtdU4ve8DUGZDK2y3A/SCs8dD+b9GRjGgy3It+HOD1v
3dshyMWk+nAmFAs849wIQGRq7Gr1f/JCimvvPF7JKsOZs+RQIjBWCdoZG/8Q9X1Q
CzxMJCPbmWD9U50paG9h2lNF947b8eNHiR2cpMEQv08Tg7PvQ1sPepCzbzrGR6dA
cR07EK4aKVvFPMX1NejZUz1tPpgx1+YamKw3j742bkT6qGdONYwSrm3DFB23UILu
UcoTqcehgmfLBFHcmIeTr5fR1/3U5+F+7HEWK5S/uhYpvNhXhD7Nf3sgHmpSMe3v
FCFizU01mZrZ4ITDzMFkF0pirlxugO6ZelqqVmhzmh7H1Qdx2IJ94KJWhu/HFQFZ
VIpTsbEgVZw3CiF2zrPb81EFj/Xf9WmHp9AZ4YpcVIVSJPvdQPzQm9JA/Ju8W5MF
Bw1DPncHeIVOfLdyDmKVVfVnfyMNIiiT2FV0xYK2kdozfnxRO7SRW8sD0PcE94Za
K5IkZiJGYJN7qE/7CnfVkbpjT2RxVaUH6+90G3y+sDQPWSJQr5AHTZzhaS550wTO
JNP3wBl12wsSSPuMkXg+S+aonma3PqpHZO6Vx03D6K9G7LPfruVKwCRRJH61Hm4A
YSAPwGVkOJutmeFwS1ro5avDniYQwsLXd8EQ+WSviFfuoyYssTxi+WpUx745HrKi
FmthRqRuZTzRu/2SU0HQ9fADWkYpa/RaL9ztA5t/JMjoreJoM/QfAdRmxRIQhQZh
iwSbY5/VzkUc28DAyGHhY3tyFiQoYkHxH6HFNB8jNuouqHzJRISI1O37iYzLAwL6
PK/Ne1c8cC+yh1HH4hOPOPaB2Fr+t3VIHKsgUB9LcpGo1gBn79MwyrhmaNOvb58G
h2D72nU0P5qb3J0YUXosxLwvDErDpfLTZHTU6UV/MByBJ9zQ08zXvki6yW5BV5eo
BUTdSdCFQdqODOtWGPm27BvppSOMqbFk6Z5Iyp75Uxg0l3aPcu9+YqOsWdmvDEtG
8u2YIpJ/Hiv/oywCZbqN564RtQu7sW/juqAK433JmVyCVUD8AC3Q2SwS5HPBd8zX
5TY3xklNiZCAbIko3CxUXrKb1NepkWgnRfkXuuPlisRcJsJn9uL2g/PsNsrsHJOO
oh0zZY5OmSfXyh0TBk4sp/8v5vSIYsunXxiPsq9VOvZYH7Kn5pZyM9GZkHWfhlq1
hoQ6hvGj26JhQwfQl2NAHdnAhvNiSUQrYgAdDlfhLoh/Frd4YgW+IQllxbB6LTes
Ju/FsLQxn5g63nUaHmHeBX+D6C6TeUce6KX3al+13PjiEtLuWHjyDSmyus4L+wox
/EaAs+/N/PBKvNVHqT4JdOdaKeibwb5IYzihex7pSm8DZUKL5rOLGwZf/1UFREfT
XIpzxjfdDqaYv7Mp8IqkhTt6HJLOgEgqTJ+Aae7EU5ZWasO/b92GadH4BPxWZGmG
JXhZyQkhTGkTQeGQXLOL0D9wwmNAh4xjBRJHpLl5HWupHkmB2d7v0MlIGVxItI20
LYBFsh+JOkWgV0VPMlkAFVIoB0YYlZoF8uHDskSnux0BbtDztvfR0cd9lN2KKzLm
RRdrwccmVBNwnxap5+JUbDHeHIXN2OLEZr/Azt3zJ6vG9xJdfSN09Kh0tvyC1CpU
9rOEbKx7S8okiKuP+NmsXZKY2C9avlv2/+rARwwpFkGZhsFHTwmsg7PYG6DWX1s4
ITW+gHU/P8vpXVOYz2aR1dTVByVYe7NivcQuNnN1zWxhS07wAM2X3ibbGW1gg1J1
Guin9gcG/3EOuiiKkLwK5B8IGno2MGAm4RylX00mMPur+3D/EFMY5DVDd+0DZJIr
Z5VwH+qXrm0c9SUszP0iiioujSSRE/m42deuTegyvGait0VvdDzvwTVHxgyHsGKi
pZ/t1Z/D2hs7SfSnzPpCjewDwK+fXDmn4zT5h//VjMZUILgw8uK6f4K6SY7DYZ7R
V/naQpLDafcq5tsgC6i6mHQNNiEdBkEjj5R2sl4HlP+bgQFPc6JLr97fyo9aa42D
2rKh1iyKVNQXYSY8xPVxZibUfXLv5EDMJ+PucqaGLifFMLO06J7ku6UJNheSaTNY
FSfAskGY8WfwIhO9K6NeBKNXGFmcNoQg6/ZsKIP6zVj4uT+5n760jlAWGfIoYaQE
RcOJ1pIYotzQmhDELD1yuhfAIuyIf2G0oU1DU6A6lojCtxQ20uH3vqHp026D/FWE
muCBOkL1jW3mHOgD2+2sg6uq/QnYEsqqbWcKNprVv6SuF0Y5YTYqQmvFWHK3DZ8k
G9BY224a1DFaysoHOAWGFgGUE6zgsy2WPGC7wMcQtj8QRNNHX5fdnYeDD6GnuBqR
/IZrAhUQv5kZHZFP/WuCIiOrNK01/25N/7sHO14G2wF/H+A0fbwQ76J1TkHBaa4V
U1RfndCVvjKlEv64VeVHe+kuXsFrnmLcmq5AC77OAdgiY1CWcj4Gl+akDqDU7AnL
z81tJflRq7f+rwdUkutDQANogHDBXw4dNSdRmnMHyQujtsjZL6BOfjcdgYtsxEVG
DGu/iQk2u9MJ06Fsf3EdRT88/3oHlaGpu13CUgiblsTPdBLw8WfyYuxDfQiawlb3
904Q77I7mCCV5F4RuCnyJILxet1ST4K4SHBSxqQ3b56jIh++/dMpJ4cRj4+g1BQL
V2B3gX5WYupbFyK22E117uE0JTEG9S23gf93awdo+BEE9oobEewcBP6WeTUjrxba
HH7/u7+r98FOa7jpa+he4eGUZwG6KsiHCTiDmWOxlxMjknHuU6VKXzSwgz4P01qZ
UQFAKRoyXrsdVkYpUR7VuQXO/ZLG5TfRc6Pa69hLqinQZZ/h2fAjfTJYmrlUClbM
Tme15sp50wIYll1uVMqmVfr2sq6W1ABzdSLAHpSnYn3dbcc+svfjjlV+FnNLwEaz
Vmr/feFrWgGoVyf8+Jm+2YAxIqAjhRiPg+Ng5Ajqqc85qybEw3DvAfUbI1Ni9cro
uqhhsCpRpmgItuaD/UK4TIxZ8MdzEM/ify2BRPyP/mg7ALaD+CK78BbZfKJ8Q/1s
3P2LoP/JA8xq5oqXl8JyOXYingaagtJKwlJ/aoyGefvhyedCk+0zUCwegUW9ybNF
DNfRNqjgQDiU3T7dnSfqjMcSg20eZfHRa29TKZW5PmU8Np6xzzp5KZD/P6hc6sJ/
N08k0AlO8wk/30e4I0eATZVC17AjtAwiIsItzznoxtVxRz3R7fdIx/RJLVkjUedX
IY1UqTyNthq0voEOvZ/3l7kVsHdaXumCzOFWfYn8ouOSazpBfi9ZRPBpowX0coH2
Vs5AZ6C5XH2fcKZa1JJnNRckryTTn9Xg4lKfMxKlbuB/tRkP46XfVbCPTYd3T7ZT
T1gmg0glZrVfflINBq7iojJAqCgZsRJrHA5nZOyEcP85AFTkW1150O0qqUrAKOCc
ooU/JyuRYMom/lGOZtSsM6j1zTpKeMZSVhlxA+JCCC0z8+wlhcADfe2g9F9vVMrx
bWlOLRJJgwp0EQ8wtnJPQ8U9SiISlDPQiO/7OcjpTNXfqz7yGan31d0bW7eVKqzJ
6wkOT3/JgjDIdWwTpQQoPbo2mgTf9LFd5txX+FDvt40J1I51GXosqtrrD08w2vdK
tJBcSub5++j1lTU1F9rxoNtZ41zpfhdZFPV9OKQZSoMB5NtVXq8Xvh4v9pc9uP/w
z0fiNqqdqdFU07CVEBe4rKmU0mYaWCWPtYnrvyZi+H4I1DAfh3q40qQVORQ4Vi9w
k7r1RoqN8IhadxG36oj2t4jdD9iM4bDbv90V3wWKtv3+fLrOsu3XrrkK+6/9JWtu
He6VXo+RDK5W9YFli6c+kixisT2RbKkxFiSjU3PzLYzI5xblWjERq95yXuK4K+1K
/MjQFZCUI80QqmiSzqHC4/BLVb+WqdG15mHBjBfvKqMG3355o+rrVNkT2tlLC1D3
fbEfJq57pzPkefysyTrRQnuPSHq8yLoU0hrQjox7wPKB+e/fg+d/7tDSKxzg9l8l
gdXrVvm1IAEqR0+lAHev2NbKb/2Zrzdcduxcy+W5JZ8eFxL0Yn+vzEpKVshMG2bt
3phAs70+58NxLLaUs0MJAQfsAMl7PiOvXMqq14hX/syvanrmBaATTUA+65uqLXw3
tSpLZOTB/BWk9TeKYfcdD6GFuhGEgJjaQ2YBDEGXaNkLdJQ8VitGi4BblyFQ3lDc
sAoDAlrMal0zuf8Ugn7nhOnkJv2vlU5UUh5SQ+8ljoqD88mrVhhnooypMi2W94DN
sEfyRPWN/shG9E2nQzEtvUNKb2J/ZchtM5VtI8glSxK8cqx+NGgzUjul1tKLPddT
9sVVm+Jq1otd8zE7DKrZw6M6Rvs3rZqM7CbflAvlwRlD6ab/mW2brD+U7pdRIMZw
kVy7rRFlHi4vGNjbj2lwr0BKC1mmi6vZD2oliyxczGk1WAufyXixaI+zuDLRAeQi
IcmAnZX4IqxLX0UcSQ/wVd6HZCSdolOa9/gm58ZCP9YW4Pa1LDcO8SRxwg5LAFqg
UclAP3oQOBps4ZnPU3SlXfFQfXeNCwCob3baagtUVr+Q/cI6YqYPASRoYkxKwgem
F+xmU09teidN9lQBwbojhu2BsKrT1686Qjk1IFCUQRSDxTJ8fc/pe6dcGyerqq+E
JoI7e/rXXCTLHl2wTq/CnH+U1xV+ZxlgNKmqQl5U0qAmx3T+ZHkvKtzcdn6A1Voz
SD1q6RYprc2dTEBLOBdxZOg+lXC0/6CfuU8R3IVKpBoeMNs8szYiGQX2ToQRJzAO
wyMtDSGWHMCtTDKgn425iiChWrVfp0QSQ+fIy4UCH5Y6vIy3YNWkg2u/zKsuraTu
PsJVq85ejYNSm7hkeijyhO7ZlS029R3KD+cuRS7p5QL/5D/WmRbrvJ3xOmChMPVn
k9tX4uoMbMeGusD3JPDOsLOOhX22BsU64l8IJbGwO1FjI2x1WZHmMdBXlilghux8
PDuVuXnFgQKRIfNQAYlJyUZ6sFQKqlAJ4YTPJrvOs2V4GM9RS1rSO2n0Gg4uZU86
LsuLLb96zFllK+ipgDIFEWxydBzM6V3xoKecuyIjT2PlTnjZe6DhmUyeW/ePpehp
M7bDuSicAGC+y/XxsFDtn8BwQ1Cr8PJpWehq5vTBLBMSdcMdud8IWCMgPSOXJ990
6gc4sbjgzHtya9Btf8BHVrAxfpxRCxu5q9qD4ZzeLz3X4z0Gbud/8Yl2zRoo0URc
49bYcYUeBRLm//+q7Wyt2Bf3ER8elV9sXHO1Imd1sVGzvq50MzTF8p/p7OJq55yb
pFNjBahNiY7Cr6YRj/6hzLRj+GmLV9/5w0KC0O3bursuXohX5EMAapTtiLbsFqpK
G6Ll0d4QdzIC7uzcTo6AlwSyxOwQxctorUCPTQb6bF5pBumKWTTAg4ygYZs1laJC
zChmJDlmGX1F4xqyk+0I3BSXIl7IgbuIXlL1Ay7YbNacb1Ek/UhmvQdhrc7DuNCg
c0uyjxeeJqO/an4I1VeJXOoVWBWmAX92IWSmtQRs12scjAW5ze09CDZnRtJWh01b
hbDSUqUzJu0L80bSKSwkGx29z6+w6B1X3sE3ZVBIpHqAmzg9L3TAtxqcYjH5QBno
m1lqex64E29uINdP8MPn/HHCUgxvH4axDBscjMFJgj+Pju2VxiMx0blfe/U3y74d
MNIyrH8r8K3XIxAiFv57ZFyggchpUpXYkxTNHV793y/N9Y8WDPE6q8eP/s0Pkrug
yhkgFJ2nG2XVHHBbBcRtLQQI8lCQnt2D5yfp4iUU3nI0vzEmtKJypJ/F5b9x6f5F
oSsDD1p1cegVNlwN84SawElVW0mglaRZWTa8zqKGdtfzp2Y6UZEDxtQn9O8AsRDF
eEYxUCS6EcC30FE06YONGko/KcEKzFswnW9jpHomjMEn/XR8rIBHkEhR1T4d70ne
9eo4J3d2QghvXbM6eTyaIoIyGOkUu42uzFwEddhTQ99f8noJmM60a33WpgkuHbMB
SEJHsqdEyTqkSUqgd+Gf7zMcSx0Uy6c/irzfUZFtD8w95QEYQDC36XRjrEjyW+FA
TsKVP95wFKWka3XISLwV373e7oLpP8t6ErYfDvOkqX7T/ZcuaNf6GH85PuKVdvX4
uzPz11eJhUo3rg6OELDqyKu8VGgr3Eq8fhWTz0YL1rEhi+umUItZ/Dri6L9zj3ct
PYQGeCwr0uhWS6U5Ggnrn9UOI2XT+Q8LyuDnPoMPtFsa9+A3LqYL/voZ+6UflcE4
0GQ/DsW3eTXuWvfy0j1wuVgmwKhmzfIIDO6CdsfcurRUQqQsqS3v83aQ2hGbKVkt
CcfK8w+SqLJZgfiaW/pmmFFawEeWQ70CxsPGM4Hu1OSFBeJAtnoupAKZlS/vrTWN
44dNty9JVV6dJUGwd8r1asC5ojvwgggKuPD9EMrWQD1zyahIN3z8agO7XZyH2X8v
dHGrBglPdChYIa2+gJb60A4vYMLVy94x+qxMj7bgP58Hfi72neEmlVTkqEbr+Qkj
HtKyRz8d/yXmdDEv0S7txE9CLWZCACWipKa5DDfXMmf83is7DLwiWsQzZZ+hOMlt
IS63p3IcF6szsSPcQHq7uOWpEFda+3N6+B40SfF9C0c1M8FZgHPEMV5QIR+a/kPI
0X8CTRowZ19+SD7/p6sxu6f8vAa/x5evUcGNYO8Ct3TnM9WHwUTdq/ajZA0I7I+t
ICtFflpEOQkjiUkWlChXiC1allP9Xo9D5HjlEHNXGL+xDXx33OLgqnVMHNO9ncZ3
9rrNsuQ9wqZnm677OPvqqMvMYXi3HSyYunbhiLjwAzw0Z77XdVM9VO+zNySQBwHD
JRtIdRFZAOYv5zNNu1DhuWIWzdq8isCSPtXS+vKPAgeOlrzeF9IOD6J0lXsx/Ef1
RrLskjN+q3wbVLWqHBvLf71l+h9f8EdWzq8Gj6K1OFteAx/sjRN4RbXoEuOgtbrs
HWPkKxXU0iUGYoSg/3tM9S+KkNOFEYYDdl7HWHxgmqhTtKy+4+yUyDefT6xNcPDe
goPtA4rGVYLjnTO+Q0SC1bJIUxDNPqfDSOCj+I8pnreezpgjvCujKNnLuzQ7ipxp
EwdOaXJci/xLgCIgPMoqYVF1sydIB4zh8OPztQApxVkqFhkV6XhH4PQxT2CKCpiQ
cLuhVkB4jkK4uHUgheXSsQepnggeWPbSHl7PVE/o1gUmDvspbZ1eOwYTg1bRvO1V
Dk5kpbjSJ0ib8i6/FXOFaX8EV11IzGGfjWv1Q+aIkN5wxg8vgI7rAJFjCzXxG/FA
HPbLCAjsB5ETs2RODtI9ropwSNJRBLTLsI0SOpYH/fkrx8i5n4tX2NM01aEmd3Dk
n5+GwK5I1k7gJknZDE0sLkKS+ZK8KYTf5eJ4CnrzlgZSOicIi8jGdUfG3uTqNbNp
mR19igz+H5z2wAuRPUPsRHu7TfCTyU6M5uL4/yvhkUGrNRYzDTztHg3DPma1xTtz
5tQo4KDOlDmOmaR1GdeQldtMzoD1vLhp3hJ9qx1Mg78biX+JS/zPfaYnIHsRdsEF
dixTsklTuwYVOgWfP7Qh8ImdgGrKXAxGuZbmlrHvx4lZS1qTI6h/wzjEyph7RGv5
LelLKsniJW7mtrcHb3sYORjKdvH+LGyngsHNX3DADTdmL3REVGld4O9rA9kkN+Cd
igWue8A3paxVLxhxKRA+Z4LVogTXpX0/aIqXXDfspUkDNmUgYZUfnqsWuWqduE/v
6lE/TeklZY4dTa8SrmY2zUs9ohmagnkhLUvVnwvjW5O3quQKqRkbDyG76NuEdu94
qt5BT5EaUyhS9TC/qomMdkKuz4Bmwk9mae3Jf2JIzCGKCtsZARFgzigRfCWZ2qaQ
1bFxb/0mTWkBD+2y2jy+P4aA7sQ+1qVugsSHN6uv+i6CePQQ2v+p9tx/fvyVQLw0
bIlXxgSWoV0mq9O5nHoYUHbMfSRyOLhvyVv9Mpxx5P43rwdtA0GqxQc+SkOPn8fM
QwuscvH6QhOMbXjvzsLv0tQZzcJFAn5R01jpARNhV2sD8i9WyEtOrYtdl4JgfaCm
jFGl8MTU9eVnjEDY0VFv3nLiDfMSxBToPUQSBcqHnqBrabZgzOE2bnMvtKEtDizb
no4FWYS7fGFQEzs7pCyOHLLQRTNv/bmSa/ZY1t92rU0o4JA+Hx2/6e/xyAezDfar
2UU+u769VGid+tGbNoYilqbdUfDIBeGFcQ4QZgRqEbqANZTJsQWU+4pfkpSNNO1L
VuCxSBd/va79E9NiU0HIaF69VqEhu8qAQbOUgQHiiheMSkXQtfZ98ZaaXqbTtP9c
YA5NsvVAG2POejxfG0MDolQWQZRrv6LhNRBGX5fgGAmL1Sh3ffXV3rAw6uXzEHt+
7Y7Q8C4+Svhwve3MGT8Y3dJiBDvDx1ajLb+HRX7XugISU48OH0RXwB2I0sS18Bdv
cw30MQMzi1AhJYOk3L3K5JOwv4Naqvi6OhLr55gJ7WHhhLXqrlD3LloJJxJt8Wp3
YIo1ABOCgYEsVCYZC4uc7LPqAc19tVSqItaRZpVt9W8dOohZNXspjOaUtNeAM6ST
dYRbbEXZkNmvCgGDfytah9JJ+YIoV6h2TQF8US/cByo9BOt21eDEP+8peLcbhntQ
AJAGWBNi/hN3rHjji6SDgURVUG0fPiIQvDWsD/qvyII+7EMzQ+rSfCBbVJ3IHQt/
LVPwgJWPaONYtdd4eUxX9nnMwSALjpUNa/3jmARjpiWUBWqfTLQjjx36h8hkMuy4
Z/4C48GKLyPuqv8XmoZSy0kEbnj7WH6jVyhwRbu+9D6teNsH+Mp3z33Sr1BykpWF
BpO0wxpQAdoIW8m8HsACmtmja89+n0BoSLdZYWsy7HVsFp8ujBHPG+R+pg0+mCnC
m1Yz4BhP2pDT+dhFBycTD8SpSJd5Ni9IMVIWkyjt+j0xWKZpfhW9NRuwB3WDaM6Z
R3bUVxM09sUJAiySSOMu1oyau/Yev5cbknJkhV3rd3y0iNgqJjBuwuiymb/CEZZV
atYNB4bgvWSNWG5XhmFrs+B4hnD9EH2HnyZ+wecVqXQBfUxyaAPDqKwwusiVyqkb
30EI0gx+84msgJS4u3uE/wPxk9kUyMKzDBSKLgy+O3bj57nZyG5empsAvSQMLLyo
j9Z9glOyl21/TaRyjfPq2ZR70VESmtNAEKgVgEDo4ML+TATXtSNiSBps7UgB2d0l
Zua4NYP8xQqZdx63hEVZqoLqPGi6dODdW8+Ccf92pUOcoBcjLZCmfPLnmNq1o0K3
K5JJmghxYeqm7USQYFU/qditCKRBFLidVBCkTiGcULc6P+C7vb9ZXvmZT2XtAMVC
n/zuWg77xScdXzPEWy231yXig9k7cShEq8oeBP7RrkHMX/0v1Pkdqi+kZu9Lx+pG
+hqbTpGnUxn+cIkzqDZDdH140VNLJX1BeKzecHrSFx5poInnd4cWIq7xvXrz54o4
CU1UHqPVtdw4Rzj11RQaEXRANST/x9cNpDpQ27kWIWsqsLzmgoQm1sgj2NXE/lWu
eDRGfEpwq/Qo0b4BhoxZV2Xx6DES97YC9P1mtb2PDHlkCzFzZ0thenTd0ZVPq6ah
IMgODw/iV1mxQ9y4C3jFesMav4RuZ6rMzD6uGMgc6aIXGHmP+DpZO/qwrh8sKoOX
pp4wd8DOEInkSNgB9UmuCRUQ2h65YKEgp5JPcxAME2zZ9Ni651N6lQgqrSfDAXHU
45zaWUM4Vs0HMaA+LFfjtcs7d8GpHDJe2xsYmAxl32j570Lf8HXyFfP4enDVEB9G
VW+/+gBZ0ng878OluZVzo0caz15XY7B2QiRJdKb6vSrFM2Wuq3Sp7bNFTZI4cNrD
wGe3tKxeUBZHWkZ2csa3YHvrCdQhtR9WfDG0DVfdLsX7KeN7iXYza6ViuDqOUqXw
oUgWUVZ8PP2JwqRDLypVgPviaoQHaSN1DFcrsJKFeHp1Mev7x82nduG/SpfYfucs
89DXZLlrSXKzqVgMrt0v0t4NlH7zJzxXzWQHrM+UBvRkJwmh5yXYJtD7sl94VWjZ
D5W/+QcYjxq6Y0RlOBO/Wai4M0Nt8k4NRfBDQXmWETd8NlRIionyKmLnMBl9k4/Q
3PtU+oOZa5xSvPPOBMmI7MFu0oxgzyYFX3AeojmeAr364q64EFybYQSOPgdoTXil
BRyNI5zEZJMKunELuLPEYeiXUs9vwiYm/FRkqk74ZF6cXouw9b572STWMj/dhEzU
Q+oWqYh3QNkHX1J+I9olA3nrvtkTPQY3rkoA1MaYFqH5zCQ1SvbxBdssJk9t6Qsy
r6ywmF4ZSMcmUpHWhp25LDU6+DWfYfhpW4Nwl/TgbXRhGlDcaCE4ql3HX6abiPHG
f4LZNOHxv01tUJaf920eyB9Ot5Him5aBtVT6QBlnrd/axh9PeG0gw0eemhNpO0ff
3lhKNn7Jue4Du3fVD6T8qLrmwap/Mw1i2eqvYtxuDKhdH+Cigrdk1yd6RBcD4pXr
pFZNUWjT67ZwwoNYfA9rBcwEfrmA0rMHNuxftjWLD8RWKGC9JDzqE3B5aSEoaMdl
QZbBq/RNH7BF8xPiLidzBfKl8jOjYHh8UIx3bJ3vdbAmvSEP6GB4xxLN1dNxJ1jJ
VEM5fBzsqg6+uiOzExlmmd7L79sY4ikJDhtJMV3b/ZNvBD/4W1myuQntxzKfnOb9
j/BqTQdlSmgK7aB8nF4xx6vWsJ7ZJz1YtNnQQDuU9thAkzH1HiQbncDiCOPW8HXH
pxWJhAdDpJUYtz46qzxZlg4Bo0YC/QTScp654aVlCt9UeDZ/wJ/Ar979JdeS6Y4j
uWJVbl5cCpfntQQPRLE+qVdRvhfB1l2y2C7DGRHbtk0TBWlQeOnZQdM7KB5lwPBr
ElwC/cT9wXqLCJaDDH9zjqVZyzNxLykHgegQGPgyG+/DJZGxudf6DeJtFrdh961K
VfLA6qQNqG9oHaazmo858mXApO6t9YI6BNNuxYVcblUIt6Ulnm0Gp3nJEZWsNHM2
yImH8UeWLIb1RLSn33wLPyCNm7NTgFp4cANpGn/zUk/XGdESIKTPEaPKm/TvX2LR
QBDxjW7v5v4TGRVd7jWehzunnc9q8YwJwnIJ8a5Au9d4WMwQ4LhyvT5YGUA/afQM
ahGJuImm1SBR8LoZIzvuHHiwHHM1ck/bX6fKcc1XSj+L4R1jxyNwoEZwN0/r6JcG
uj0c+z/NvVjhTLRpwxmAM0xwByR15tDg3lnXsk4IK5oBDysoysGhY5h3QaLp7PwP
TuEf65sbvWzufPz9+KqEvkAKRB4nU8RyX919gIjsxIWGbEFE8RoxsyLoJ2uvbHhK
IB0m3ZKBT9+c4rVvn4ilPGoSUvLtDteyYTSg3Yulp4i2P8DNPasFs/EELV/aVfW5
tletbpfV68No10y8CyE3+cLOrEQ03c3gnFISLRijfr1oVUgauIQ8ka583dUpBnEq
8B9Dq77ggKgQzTi8tPFuBBanmhnGNPhOWGL88JDb9TzFzm/ElUqTSbwLErfBXay4
93ADa2ygdxQlFfPJ4WtCEFDWV8/akdEK8wrI9WadjrQBy7w8zYz5+3vXkWVsvFs4
G4CMmO26cqc4Jc13Rt8Y0URrX+IJboIpjpBXP0yP+UWu7a5Y99dUcScMIPnWYwoy
g9cU5gUAre06d7i4ocuMieu9rAG3v2QSslbqBJUsstDVTvt2urUedYJNyWAzojoz
Y8kaQBqSNrfG+XgYw4ad4y9I/4R8XenphI2+1e5W0jY49DgZ0Np/KXb0bb3h3k/n
qI2WXU+2Hq5HuTCNMjK58gdMAyVqLOJ4pZQK9aZj6CPbeEt1/92Zb/tpJUyerBMY
1NDiQMIjwhhBbOeLVYA7LXbumztrxj8ZdFA/x48zHB9RgPAwQw73v2ZUBpt4geI7
1QuLn+BiwPo9pCJeWad92qEBB4S+QyZyRI/39Gfkr3QqLgupwDXcB9hQr+o0sg/T
yrDBgWmh8/pb7skA43OYlPGfzE8U7MqbWL3KauKk+SSOaknFxwU02xxWONdQNJKd
ocQUbW4EuRhd9KrEx23WSfx5fGlJwG+t0117GppwASacjb/Mqs5JSpzTmNku/UW+
RyS61xc8a3XuniQk1DuB/wzps7oagnlfvc2SB2jE6lW8sDrvH0/sz2DY4gr4Dn0r
0+0lO+0dkOo2efsLNi7oVZ07m4DD1f5H2VsUByNnrrID4NFnYj5icxe0BZhHciTS
z1wQpqu+GTFq+T4VVA+abXY1MEXmpbILYkuTlAD5KffGuw1E8FIqZpKg9ViCErSg
YDPl0Qr3TCVeJI7bakRqEEMLBJqLEnJfEtGJNyiL8Y3SECQsOxtYT2WcdTIidFO6
NHgIGcEp3NZOlHrOFMsw5IIfvV4ItPvP1T8DHXX//C3VvX0s2jQe0XeZ7jDgB9bK
6J52qpKtTynWyfrYFNH9NZhWBRX8fGiiFZz4eYRBGBDaN/oZ6K6EGbY+Bojb8joh
qdnWCv4pZnpFLAy0N3f35KlPCayZlKVo7f3KiUz4mlH2F5KWPnHTK+DOAdfR/X3E
82I0Yrz74Ec9CtVYhBEP3mx4sb6KVZaBhlKL6f7V8YbYjSVT/5qnkn+7uDBRBWEL
ZPGD3GkliIRdHoDFlfP6NeX66oaUkT5P+mu9lBXnyEgDyRwEfgT66iHXXqCAwYhq
4pB66WIBhT+ofkN/YY++udtAX0WT8n0prstfwGKHKlhVQGn8mWbvo9oha1mVRO9P
a47Kkgut8XDlr+mwSo1NDS3MsYBZ+615jgS6z+f6GlN3n76z6HDB8E7/y2g3DozP
f2Yy8xRo9M8X5DxRQmWhBfLKqQOKt6WQIAPdiKNXlWz4tVzkZ2fx2CZ9Gzf8i3BK
UoH9S6DVAtsfT0traxBTp/kARRvTBq3QYXDF3PRAB2DUCoAkuEseNRhqGOb162rI
cG69XADhpPbZoXtXLOEmR7y8GQgDYyinfwICquuu2nSQle5luA480NuhnFHiFffP
uQs7+eZMDT9/OlgcOiDh4/6ib1U+v652oyIIcFXi/mRlQd2FrkNrOCCaFNfA0Gvj
Eogo3yWpBvqPNdj0wOsmlKRiHPyVIWzO3DAgovGsMKWYbVpthXYyAeVQv5dyRBe9
ucj7NMx+ra0CljaZbW9F4E2O5PQe9ciV+/FT9RNNL7z4KU6sxqPAdLZBS19IddJG
2e/ELi2sxuJPPjoWgeO7fAgw+TVAY77tTXGNh0ayHmNtTBTKr5BkLZQ4c+BMLPh+
ynyAoESWTSbxXUTKZ433TMK7uU9Caf9PLi7nN6u5kc1Hd6LMjKB/0+hNIb/Mdxch
AeY/erpWRntYZiKjhnvI51GEGkEMbXqcAfTOiREBoQbhKRjHBHJKc8CPWKIELnE3
+0ZyogmzI935ibJRGWUyke2iGjNtXo0WCw+mG6BDiusrozqOqWqi9oae/pIZkRf6
M9qw7g2rbc0UZkByQHM7zr5IldflQ1XYcDLmTUVVDOPD0ro3lb031ztRmsAoIjiR
PeKgLzaXNlXdhVddjhHHIpb/MSRwEm4rxkj92e45Fm5vgH7iDRGWOZRJ7f3Cnx+z
38UgmckpmADO4uyg5kh/GfMKl0yQ7ycEHYzFC7KHB2iZ5FKCGdr4T6yXBI/phYgC
vf4PXWhp1Wiw01VuzcJitJgegCf01ekdJN0M32On7pPqXDi6wXzivTfyVNBpTzj8
eWxneVHHLsDP7I7dory6zgSqHyQZ2TCYh7z5EnZRuT+pCDp3gExBwboNFUYGvtPY
3HfLd+pzEVpSqWY3ngHUVTdFbhy42KsPodmesKT3BeQKp6zfkYyuSvwTGVavLItE
cxPvc/chY8ef8ujAY3fcCeXKubOmq6oPkVFu95Y1AW537wG37/N2zoU69WFxhf4u
PyKgUZJbDFUCa/Srq6tKi3fsR8lBWErb3rzGgykpCnVm3uF3OD08gTP7NTENxKk+
4hO3QLvKKGLtSxYgBe8JyzdQmDBGl5pHhTTiDhuhz3cwphtDYomLujnzfJTL94QZ
qjKM58hF6k6DWNAf/O6sHm6ArloN73Lb95N8abPS9M7cngq19gqItRBBClaxUCZ8
vcwbwSluDiPgFNBc3GgHvkc8e8gtf69ITDKrCX9LYzIcxSBOB3xsupBHhMEMYw5a
8XPF4MJ/sRzHceZRt2mgrPOcA9NpgAOOdnBCuB2zkSyQCE1AggI1MgcRcZgIOq8k
ZDZoKLFLKTzMlxN0a7AnYAazjTkgyBDoNoARO9GmS2IdBA8UP5E+yakLjdL3ngom
Bbv220g1+yiILK+CByx97UlkmnVSasgvU7d67J5A7lv7PJ02BoHSLc0nJQNZLtKh
YfbrXtEfIvBKrGQmntmoqDbAt6elua1zBB8yr9yVSQzzJcaABnQ/BQ9cUEupKwW2
n590oktBwD3yDltN1Cr5JK3au34NOCfDlqUULWAj+Ftc5hK/8XqkQBAhHk6gvKhK
C6pJppXkc8Pn5Aynh9/T5rRTdt1e8IA3DZ1EKOPRpBEIAupZKQxmU3mCPrM+ta4n
VTKaM/Uc65zZNVuepxydxen/taDm7V6SfRoMG8DComs1Ch3h9Aaxlzav24erkYbi
eoEvJgm2swhkFqkIDyj7a989HfseWHmqEfX2OsLeQiIacRJ5JziA/vizmrs61s5J
3u3jX0U6znbuPWaEFPWIqs/HvYuAlNKKNhAka4mO+fmxLaapMloWqCPszvgznTk+
qfnuEoCE17VZhw7Wkfd+3PbbxKQVrbrhQZqqy6EO4hWezgfeJyxQW30MkLkokgLL
bCkEghDjBrkgaQ7oy/q3R2/ALQkc/b2WcRj1BR8gEmksvP51iIlZYbnWx4LiWBks
wD352ShzjEn75WSxV3FUanGX9DnUhQSBQ1iubYq+7GnhWvXcUydG0aQtGSMCbdgD
9bWrYVm8DfZsXTeXAi8I2OlKlNQR9qT5avyt1BNIF6b6U+8+Ve/KIIWMBR1M9tht
exxEm6Vrikxhx30bdZKQqOOPDrb9o75CceZ7WKBE/wAS/+o/u586wXrOPBDBlEpy
t8WpjxpDW7AeHeuiwIGqW55iGDAqmzelRXNTGwQMQmlQI6FkEz1T6JQpVubbj7HT
o9lx7Vg0gzvc0kQQ9bl/zL13/MFSVoLf5k0i3zxxVU6fedSNyH6yOjRpsCcmlGXD
tvZMU7tVrwZObFc1W1pbuDishTK76ulFxbSsrxiyXhPM/meGIEej1/9YlMWI4UsA
oSnSNue2b6qslbqgJXpLL1v0t0fw39wLUVMD/pdMPapJ8NObDbl2QhMxkHlnsrDa
d9jQDrTxCrJvWxu6uMJJivbjwA7Off36vT4icx/QuBCpSmgpnF5zcv3bSEQeeX4I
vYtDxMC1KdT9V25vDz2zNJshd0E38aFYv0l+nr4dIS7cCJrqQmUdOA8zmn79gn7u
8BpSMq8ahOscVrjsK2LTZoRDUvwXXxZZAdMSoU9gCwLNWXg8SrXwFQFTAIRCK3MB
4y5LDWgQQxgGHTKTHBMdqRqKR4frCs+kltqPFGmk4tRmO8+a9S3whSqYKDgtO1sW
+arjBapCXJwEQBFZyv8WwAwbb1CY+ta9Xut2ehM3qvchwiFZiOxih1KrZzXvZw3T
LM1fwVYJH+hHKxrJWZynLGg0UZwsSKzOUfH8t/KSjaropK4Bb+uqdUXvsg2djN6K
Q5FMvRX6ldfPO36NYM6FVNhbRtlTVidK4+5fYG4ZyVGTbdxkRjZsFIIVusIuBDn/
Ic0WQngNNmmBOS7JNVpIPpkH6nQPIOh2cqXMKBEpxDc9ZdY0yNkelHK/pQXQwbDt
qixqfiZsksIY9I2dm2U6E3KqKUfpEqForBYVGnQtFyL8U14oSAIZ+nO1JIzGA0Fz
rMAjG9NYigaE73b6oFx5mBaOBg/mi07s+1fkDLgQG9TA6+PlwTi02XM6KeEBcRmR
3WirrxMBldEjJNIf2KsSszAiFRZITrN30BtJc+83AQIl+kvFk4rnR2hc+F3lh0Sa
hd+fB2CIzKkdf6du44n5C0z2PdYywWNle2tnilDItDWY6T+uviEFzi3o1zxnQmpo
nuayTQxWYdcQxwpUs4oFZidXdH80+P8whV7g8abEUvHNac9llhAthoLH6MuhAvpm
i/TfEVww0lWaW4+6duvUptqaMgrD657OAtQyVP6q7xsoaUTaK1hEF8VCn5Nz5aRP
ha95anmL/rwco7A+u+sZgxx6wi4dZ2W0nIGKn9dM39abwmRG6LKE+0ULkmul4hVH
r3jYah4NOs2347keMZfoqZkvgVH9pPJwmXpwmha48EJw+f4m+Sq/nsGC2JRalek6
Ofp/28gw2U1q4mI70hZUK0uiApzZ2lr/2zCt7G6CldRqO3lEhb05mym8vQzD6FrK
Aim3dXMApwy9wpY88umCGPTzP9zYBiHMXnvBJi7P0q7zNxEdY6ryRwX3PyUE3VDf
nCnGXTN5O8ButseP2ychRbCZytoTF1PihrN2MVoGeEuFdNeWFh2VK4ub+cOByZKN
XOIBO/mmxtxWxgCMIVKOEAKskpqka/jQP4JXyNdS22902cyqc0cmHfq4njpV3WX+
to6MAkd0TJZHssxevxBn+3Uvj5PUK5qCHO8lrdDX4CX3hFOAu9pCoi5bkuQcs8BT
5hEodAKgWrm30eg6nZU21GvBQAho4kmIrVq1GYdfDlVXiQQI9Jc9JM6OCQLjwCH+
yASQS0kAsxQgkOxuKONleSTwZQn2sqINug7yrjLOP3EPnu+tyYN3bbnFwEkLbZBO
1hO6d7PNXriURTJygSnKvtbSQEAkQRyaVKeYT2UkvrFYAtYjbxOBPDzQS74Fmko+
SFWW95B8cCUMqNyHpl5DYTJyYqMfOqYtsSIeUDzFPGlyawJQi0rUN/MWMABMJNuu
28nJuFXJu1QBKGoXj96kM1TSsgONnzsg+XPQeivJINWImHT/F3JYLmYjHWaA7qW6
cnl7TcM5Z/eJ10qpl9YkaaJVY7SLeoimsHfPiyqkZOryv+URAc1ZK+VEGifBVcZ0
cIZhMMfj/lLo92HyIUA2Sh9jHiTgg96tsCfaBjD2tOycV2q5kd0ugF/4d0umRBX5
+s9UCdht0UaKMfNb+AVWYtPGEDvxYOe4U7dV7vkLs17aF9Kiazwiyj7aVwT84Bh9
tu9bE54M+tBfaVlzARZ4XBus9Af2U1z28E/bU+XgknlQMg82hkcB9yNtCYkrHeFF
KQ/u8RXvNbpPGXOQD+TXe9inYZ4YM3XdhSNh3iKWLBIGXAbRtmLgm3t+jCZtQvg4
v6RUcva7+hJqqk26/HE7gPv9l3hdMcFPOyFS/C3KdVb1jkL+jhzBl2pkJ7DVZNzb
XBOs3p9u1xvquaksLIRTtBvutD5o2ow23NwK1ABISnENnp5FPea1AGxztAD9wXOe
4Fq+0lKedFKp5l20glbaXS+8dKfyx4bXEKW+InCLbAM9NwKAnuNE1tswkDFBx29n
91MZKyaGMbbf1HDkpOcWTao4PLdCIaVIZTYzBhPlFoshtfaAU3Ixps2xVwziEpe+
EQNaLdD0sUA3GNs1/4TSz1If5muvmnrcQvC+dYvBG/+0vTrynUJrfmRUf1hZzqjj
EEZG1EPrO/vLOIq6oZHjY0eqP1F7M0LoCzG/kbUUcPixtmTYMHo1pnHRHxZT90O5
0zrVPnek+wvuHlmetMPOCGqRYWJFNpyHMnUPrTBg6U3cWT2XWY8dkZXuW0Vk25Wj
dIhepHV4ncDNqtso4QFVwa9DRmZIM4KRJ7+7yv1gwSeMgioAU/qzLB11Vrgrk2xA
wjqFcKWOmW5uJ4zMvKcXCiWLev7ITtROl1NsEN2fIVqWe41Hs548Ouxdr4fV7VMH
xlITFlrPJHJzvsL+QSQQ+YymitN7SoK7hFMIYyWCI4DBbqar9WSymUSEpTdlw8rs
zQXiQMbXLJ3ftSQ50wQO9JyAovTrU+Ljp5s4Jms8MkFwmzIbVsJpkbNI8qTisXma
Lwftba3tR/RXAa9N+VKkVy/wMsiwTIL5Iw/+LjAPF9GnJCXbDQgQTNC9S0PuwdC+
laIaOnfDBWcZ9T8fkZ4DDVXrndpMGyNPTeLGrfCTTkelD08/C+WXnc/GRwGF7D/h
pVHQW050i+xLLr9WmFYJFOu2Gcaqo/POFPziAB7lmbOlpyV0kqCkOkfG+FdTU15C
Om3/rDSCkORpvVYEAxqFPkIxg7+14NMish8swJ6YTu4bbSo4xLmPceptz80X7nCh
/YLY0IiRhzI0BoFeoTHnLNyi5N5lavcrriudL8hPwNLF2fB1mpzMDCL0UfzRsUN4
TerEJ2NBcGbyEWu3NuzO2VeRRVNT7u0cY+2NQHfssHd64ARiS3q0emPk5J6ldgxZ
k8Sxu961IeVPUtUYBWKjuydvVDvEM6aBONt1NfAD/r3cepQH1E14RukEn4oymiie
NCPAWWARM4Bqv2r+WOBHjtclWuOcr9htGACvJ7j1uMPsdoonfwA5Nm9hdE33hiDN
TlmbhhvEVWKA82qS9RNNwcjadp8douHi6eLAme1y7j51ea9+/IbZxp0xTu2o0h6J
OW9vFQ8KqCRW+WoPiZ3S33Cgvi1MKXrRrvPALPoFJRYsDDQrvW7GPf4nNHKpeEwM
xKaOssjgS9RjtaTCoHaJVi4LXYCJRulmonYFAhem1Pm62En5pr0CZcxDKkUR1pdo
LjFbbEjE4lk4lqmS5v1gwziRR+iFEUBVgRbd5sSJGKjwMfzeiLG/zjtt/+8IQKl8
lujRV41KKBZFVKJN5HBTdpZjZYcV5ri2QY48i9J3mrcqJ75EzcPEa4ONVZWmCFF+
W+BBKiPG4vcqF5bvkiJkm6R0zFvmn2gtPT4eNcrtWoumrPNCWByBHldm3egZSP2Z
VIzxLZ0ufMY0mJASLz7LpT8HaUbli/clNuaYY6OUt7TZplMOXxLXvvpQzDcPjVze
UEg+BxNMzCt2Hp5NcIHHBU7tHSTuHq3O/K6GcC0OlxDPSYbsmBD7O90HLAAnqeqZ
HVwwmsfZGnmZBYoJhGa4ObUI/7tYLERBaLndG0Choa9bcM/X5d1CMWTy1U33QK1h
WUdjFQ+3JW88ShV+jZ8cQ/TkH6AOq+4/9Gzzs06KLvf01k3g0ScDcyPCJQvRXm54
e9GzILDIO09Kw8qEWKccJJwuA9pKz2ws567dpfBpSjgD3sDseVhCBpVNPM67uBKP
oTQoh6dTulBhhq/3iZDMSN+Eip3aFy/et8yccDbwK+G2V1xPvV+KW5J0igCfGqOP
HINkCHFXEh/vZcUDAPp7sQr+wnO0M4TFtbcoFSJESgGnys9IqTMcVRdGdrvOvakR
yYyO3aTvDuFFkblgb4oRTnQgpJT2GWPwtl1Ug3QN/hkNfLE8ds8OsjDoMIRG+X3j
qSbFsYQHHMvEH2oozA5JGkY1ooGfUluBH1pFoHcoea07614kjrbt1QAsxIl6BK96
nijMojU+nTJc5iymBp5dmrBKU+xC73TtAnzFgUeJLbSXG+6Oyca64vxUIgDYOawi
mgcMYXsIcuCRurg1izTxxHx3h1t7eqi8QHeU76aVRySfJkYGvYslBHID0AVe2+Fe
0x0+EQLRP+wlyC4uw9aBTs2/dBXD6Lik510JxwkqNBZpqdLGZ1omXxDDu6CIBDJV
nEQzpkaiPEBZA8OG3Pk1IvGXY4eRBCszbTie47otpRKuiDP+BPNWJStB4oBBReWc
8H5v8fiktQnas4uldpAb1fWmcCWPke/DZgUe8bIDs6KIal9koK4rbcAN3YFwrl1G
l8rhb7Jktx/dbt8Lbx3z/JCbeuWQY/mfHk39h/0paiChREiusHIlpPgNL0EDwMOD
WcvB789kAeaILx6Azf2I4KLXh0/9/T+Akx9s8t9yBviw33xtq5Mp4A0TvcwkchyS
AcAB9v6zJEGMVOr5U9lzdlSRaqKIH6fyer/1xYPERvthrc+zmNYK8KeM98EKOcJf
GHWznIBvDMcnzogkUW+qDkaAPfnhYkw03zgyjy4mgs3eOIyIG2McbarRgUgdBM5l
ye1V0fgDB2n9p0W8DqYAooID2FUwrzAw15TJ6vAds96dX2D1FrISspOCHjUwRlmp
RliMRvhLiN5Vt9xk4aEyRzCvwDNf9ZUjKxYzj1lY+NwTtjaXAq8XP45NfpCPIrec
K7pUrqzETLOeaCIbN9kwPbgHxa6KUwEzChxAqcbkgUlORg3lydL54pweL7F+MWor
P5JWUShBtZMIcN1Y8DDubwVGl3AVKvOC6bOB/QXpLYdQOmsqIzJ4QTHsWNW7TkES
T96KtGZA0KFNEjhjATUihIcXe7/FveMXtnwcq0cO925sSTwpKWJA3xgmvwNGGr2b
pUadGk0nHyeq2As+xmiwtttYzwEyEQI0SnmwHHTTk29OFzhS677vKtc3dMWH9aDu
8kg37wupQekGLU06H8zS+LN7dnB+Cql3RjNKn3Sj6a0jUeffs8mZ2FKjMJ8BdNj3
Gv/AUt7qP39qTViLVhgL+5ZAhOQ1NF3lLd2riSHrqnXWUOtYa88tz72WU9aT8Lpg
rZhvb1ZgUX1U8ms/Wzsyh0zsdrOvJ4OfyKO7es78oUwljvr1JcfTvSa70vCensfx
wicbShVR+QFti8ySJ1fJLBa892JLEuAZWmO10QUcH+1B5ZvOweW2e7WfZW9S4M+m
gkfrLRk5QUbwPgRMTd1dseDmdQhoDdBWxOz1hm1eglfQxyH1JZNSCC8hp9GPSekC
sJQZtToi48+NGArV2Tas64/8Shl0pMLsVpU/phSvKBZxBXo34ZzFKNkuxygiMlmO
XP9Dkd1UKScV6JeAqRmUwbuFFWh1SDDsabVRjd55Om0HKOK74FAR7yuUj2zRUb5c
BDLA+Yj5RC4g0/LMAd5OulUi+qeOaThYqpwL9XRxb/Ga33zzO5ny3RpNvJn0OZ2J
0ebyiEf6i7DkGitBrmRQPu45S9R0cNXPdMqXsVdRdbaBCy32y2C78mcPcP4ie9GT
dS8b3NTvDrxQzqT/S93W5Qd+QCShPK1EygvrOsxvUshBAFfNNLVyezbe38H1JzaR
a+SMIlVSQ9pBMrIbFACU6MN0Riplf3cp1vzhxSAHefEVAuwW+5zd3jv4IHr40peS
qKjHn11NK7USHcFqTR0EDPkJwhk1MLttyNCinm8P6LY4V8CK5Kn2h5jZKL2pMQVN
QSZ33JCO97MwomFJSUFfaWmWtfFFynRRnzlg3sRRGueGb9u8NPZI32Hd5rXSCvwd
oJ8nbg/m7VIt1GwtZ+us3zAkFNEJ9+H0SUsHcFtGKDbBHv48LxA9UnkumjuN9du0
z/XtEGt/TDAVYmKg1o+4Kz3ufUH2XMTHeoDcRohtdXb59jzl8vkLNBZpSizTWj+5
DVqoWI94DZa7TvfHb+LVY+Jvp4mBBV8XXjbVbXacRKP+WNvqKeDdEm1EWe67zrAY
YNpYLr0JsHOa98T33QGj2LFlrlMnV+BVjhMi5zysFPMXOdK/kq5nhAUtgMF11k3h
DZhDQfPlZ94WbR8ZGlzKZbw1ULm6Z08NHhXXX/5Rrqywc/BMO+ytPtvpuTTc5sVd
KgEIFLg5lfMfcfaTsQO604BtgnspUaSMnLXLEQlc8Hh6+FTcR4bgbxXLqhwiJ3MK
LMD/Aau1B6+bUAoMw9KZTknPLm8HvW6N6Ss47N7wD4zJSCIRnfiCTkZpo6MRI0HE
yA3JpW8kzx0d7fJdZshIAaQk0PDbVQQaiKbCxi0RUchR5Ca9rnPAxW4z/54vK7zj
tg+S94L+oKiwJuatUbXrRWPzpzWfhyUqwpug3ULBlKDhGFaB2304OtKCN2IME1Qy
q+bi8B4Pc1WdmOKIw2XLrAsU06NnAUJ+qboSD+EB8AVUoN+qS4RdgRs2otQ/l3M7
a6ZW6pHpbEmyCHpyei676XA7WVRqIv9nGLGL3L5RhSh+2pbJMThQTQqamVkjCrVt
3gZQgTybVwLz04Sl6dQMgmfRanrCr701lcwvv02VJzw9iNHwbqYXG45qytoRwYKN
MCvWAbyjr9TdXatmntrwVuKvalIRmRlRHPvG002tAX+EngMcglUP+tRjHpObcOYl
tyETf1SV9P76T60MEbdDQMyLJS7bIO0BtwQ532Kd6uMjixpx+HfPT/umhuxmxGoW
cG8WCi+rCjBiccypMlmTJn1Kc28dj5JGnckEhY27JvlquxNw8vqupInr4s1/RoCD
zYgLNlHlYg/Ln3uLU4Ki1HxxCFKAtDFrFxqYsXaq1hGpdaTB48F7WPxGauChNaWv
Pj/yuVR9U+F+6zXmfF0jzWVq9QCGb00rd1pZ8EaReEIDHjQKrNPvwJhhOd5n1ASx
xRma4H+O1QgGZyaxTBKy9b2AsGm7WkLvd0ccJr+A0lWqoZUdNqTlW55Zp37BLkd0
vctqCYyvkhOyohkkRH2wDzNTB5/KfWbHIRPxiJI2bf347vHqvLZmL8UJ2WR6GSqi
SrKbjqoBh+tD1zC4zzgzP2rIQ4Ilf3oW2jkR9WLv3gmouWjBDr3ZlMBNoSoSkwWw
MAr8EmJbE38ZwHBccWDXo77H/+90i5ttHfkFN32tgWjHQWHD9rqSU9HyuQ3sIKel
Olgm/ug2BYzArNENYxmm8BvLz8aPFKix10o2HvhWQG0bpdDb5Lyp/tnPEEezTITf
PsmL7TeeoWDvvfNSau0+mZMO6Ri14DlTJIQsk+jyGXBHsatmt2CXFpg30ksbEzQR
A36WQQzNhHAfWEcygmsOWCpdjX3kUr1NmuY4TXL+fLCM6El7Daiv2kb2ZeEgykah
rhtZZsoLCk2dqDM+z87Pbz3E9c8ByBceafaWB/RcNfdZMvhoMR0Jusy4/C6GHB0F
VOPFcH2uBRBFsebUBofwX1oLkrtfBZLssJp6tr8urFfm8N6Tk3L67i8wtt1hOBBG
SLOFKBBnu6QnUVp18fAczP4IqCs4yD2A8NUo6wpcEV71etkzUJSpFkf+4LPK6lRs
l8jYTcVEddUmE7Vy7HTvDDZeiX/bYJH/6o/UlwuPIfmTZ++cw6W1B6rcFZ5/dftT
yZ0fX+IvDV2tc0AKrjVXDi5atII4wB+aJGQHwsmyF8Xg8WvUm8NbOPRwRRpsEqFg
kO9oegPAtqjV3KjgMB51SoLVTDuPR9sR7jtTEBJg96vPayIoNYGFs/g3cc0IQfW5
HYhDavRS2yyaHXXAlqqxTDWuY3v8UyWqvTpye3HelZiz+9Uz7wLWVG2JL/g0d/dG
VncLlnevKvtuCs5JBq4Wm+iulyuaZFNNVumHy9xLbut9sAlepcIDKZWlIcVvxya9
lRsoiBsGZlqbEXC+VcO5z/qMZ86LHwMaTYquL7xxhGtzjjTjYajYe9CIPxOlNGj+
s/gvZA49D+t023JfKli5Zl+d34/CeRjFk/Ub95zPfNh7ZykyzMIhao541Ul3BgSv
Eu1TODDex2DRxaww9RxCtD9dul1ObqkHzasDA1uMdvVdxX7V08Is5GeokM1nCcQd
JF9YrUvu+vQu6S36sykweI5H9cffBp1LhG/Tw8jqR+l7OGcFAzQiiqnlnFPrpOYi
gHbQsKPtBEyyMuErsjzWYM1CYzKdqb/ieOI+o+wdwQOrtO6MVc8HCKVxDnEkYLVv
M15YCcaM/1kGysusZMvzYS3a4zv0TggkPXWyfmhFE6o/3Au/ime7qcRqTslNHoax
gGrFr6zlgRMqJBoFxq8InduBCDoWilJ+X2qbydafK1W33YfbVJMhVYBnKkOXzjH/
1ytXHnFwRj026854O8FbJzJbf/Nb137ChhnH5RXTlpOb+4Tetic6uiaAdAnA8dCO
YeHpnfmKepSZUBQZkchJ3YhtyKh+FGYhOMbDdftzGy4dItEkSk4QlA5WoNFC8Bsf
G6LCf7rtiYB/3RQl0za61UETviwSqhKpWQESBWQJyJMobq2WBbXdsEZoqCwYITa0
zwijvWAVMD0WQMnr6MAr+CdV4VBhm+ljmlcr826Nlbb1xqNVHO/E9bimJXAKLG9m
N2zh5djIQrOVDaWi210A3BxZhUuILO7Bvmk5va4x1D6GQSxPIvzPGi4KyqIdTYXA
Fv8UYpH3fCMJBStHGi3SXVCUiyjdD1A5KUnUAvKydBH3JR6HOAI17eXQ2Edk3xYq
f4Gs+QmiVau7YD7uWo8H7VfWDks/CA+yxnBNfSdur8x2WS0/7+daH5b60sLSBGDK
650LVKLhXKAhm9i91r++s6Ay4VYknpFarnsLGiZAkT5uHM2G04klOYIBo8R9+Jzu
y4Et0OYXGRrrnipzFoEo4WTrUcJwiyEpQLd5stqRchRNUlUK7K1ffwOlrICnZLJm
lL8+NdSJjZ7xryAoSsAKp63Uncc2sjh5ZEFTqI6IHWQyk2GGEBAyiZKzZqL9MyHQ
9kTYS2yQ+PkCjmPM/pVlzoVEKxFrnEG4mcEpN4L8SIyeMtav3q3/DpPGr0hPo19a
d91HHrKX78AlIv60JDUO7wkkSQVWNs4y0BTzm9T9+G2sjUkgOtcV5G5RbLLANpA3
xWbEAjFvN10obEXZd+rA09AmZqaravAwZxHll8WDLpHL29rZXVXGplw3+mmYta73
cVUK5Q6PRrBPnbe4A65RHYeQ6qp13SuuuTl2NABgrRZmxCTyhTtGCBr8TM7NHyMn
wl8giJ5TqH+zhGP7tcj52wsMKSb+2NzMBYNkHVJjzt+/LLGoXbZF6ojhrAi819mf
k2DU2fas0pnREEw7c4d9zgOHfGY8k+N5Uf3Bxbyoft4OTvFSRbZbwfU6kF1cDyQt
MP6hbZK3aylWxsKUzc2o1M1kkMHpO4HZlWzs1FGOFTd/+N5aeHVPxtu6yhtvmrbI
ALOcX7DbjJJLv4QzSj7LGMVZsgHj+bvLPXvOQECfGwxPWAr0y/PeloEjYcHRMtKm
T9ILYbeNyL5q5JJ0Uf5ta5o2cg2k+u4gLuQLno7A0Yziz+39m85DkXazdO1aIY1P
mi+gUep9x4Op0lhT8xfU7aGeQJCmbXsIIWmw44h+hYdwohGOqep5bOK/UtNLxPI+
FfyCRZDOHXkBk9xYKyGTACPZmT7ky7McyUTRMlt9QCzgCXxmZQ2G0hV3IpCfx5f3
wlm0a7w8uC5GXfqhaPACjVAuNMyIefeVKrSxcMnARxIEhrBWViUL5RCdcaq0kJ1D
Jv+0O+/SKNOjvrDrsDUD0EavDZP6IwMqXaUO/KIPSzrJVLspW6Dt7WMY0iusWAzO
+sa3C5De3m44V39qNgExIxTHANo+Cr2EwrPhxVPe8HUOT7pApLBM4d6x9y2mjHBR
1H4FAwueNQOFasOCMATJDx+tJFvBwCf3M55tDwlRbPDEYbXjRX33Atjc3l/+mXyg
zNyET/uSG02GjQyTTHOzCRUfa+3X7G0251A8faivKYjXpQLaQ5p0B17tserjGM0n
612QDIRyk5CtvJwP4gkYM871kRyXIh3JqFzHMLc1UM/N0lzD4rBLyp01z3kv/xza
RoNRiCBAfaTPDU+BJOkMMs9jQnZItxBJL9s1oKPPX5K1+cfK5QxkjI3aEPtMl6ux
Or7vNv5F9mnLddGKngKzIc2xBdBXsc6nxOgq7VzNab31woPYwjDC+6+9+eLGkVbn
c/DJj7FpNvaHsyRXcCwmMJWc3a5ZX5qyVqxbpObmk/iGCpD6EAxBR4JlWtSUbYGw
YCq+C7QDJu/wmtiyxrEs9hHHOR3VHZPFQLNbOvChtiNk+/9VJnKnw/v7mVK1xXWo
r6v8HrJevloqs6M+l/l2oVt2V2ToR4JEqN/+6R649m+JR6h/32dkd9lSutHxYRzX
JXthbxInTHEA3RBEBHm/H8AJ6SG24Eu/tbBq/3e+pYX3KBBWkXTS+FhxSpY2PETV
J18JGORZS8LWvsiG781RR/gWl/4UMYt9bLro/nXsJC3IHt3fVArYPU8kgGP+SPuG
wyN+FGLa6cj2a4o4wFM+afFUVa8PPjTX18u88Ceu2FaLOA5ijooJYAeq316iyc8Y
k+RJaIH5c+QAa+FiiJHGIvllAmefKDn13gVxHElNiZNxtDyZ0Rt+dovu3e55l+Ky
DWOmdKwiz1Ms0laoYL5XtBeuBvQO78s+fOw1P4jp2WlzCQzBm/MCkDGwlUUvsmUg
oDAtMMReiyp+m8vkRoaq65lUVDnIV0Q9q3JXF+Kt2wXvVF7ny/u3Jnj46FfQCeP3
cmmVULF3VopJX3vHmZ1pnaEAgdww1QtCRxw/wGWfr8Q4X/qoP5o85CEPDy2KRld1
/o+fdJD8/E3CL+SVkdhRJo7AlkGBj2moSxCs6Kgm141qcewUusxpcm5tbTJnBTTC
7fISHKmcaGrD/rMSrgKc+OOteGl+kN+hdk9vxO8oao0Q0XKifMbGTl6bp53efCyz
mbaMkAcWKyP0em8N0bZFO2G6XEp7z+oY5GPAfFL4gxtBiPUKXL3D85McNeO8KSTf
kVYoCFhRV3erNjrbiH8ulNSMP0TXqiy4eolS6tIa1WOifF3QuXkUXcCNVQudMc3r
ddk/12w8TxjPiT4hIzGT0CkfmTZndmmj3HUScedHhN5oksLQTNOnAt3iyuvXG7DW
6yOvBdPqzkc076pL181AfDXyCORO15jI5UImfkw8Q40Pe+tZfHHSsufJ/+GTW1AL
Rckmjaj+sVGAzHFeL4qN4EDnEPETiLwiS/pVF+HzQFnkJW0a16gb4GANQmoDdQqP
jcCNCiJtBvs5AWHcWbqSlOd6qGmtesF6VdALFX4b2CUQIMtY65out267Bh7Kraxc
dVp84312z46j15b3FAi0SIKMSSlKrUSC4TfSQFQifIc7vxUtl7NOgUf5AbgH5F5w
UGgHlC4CHEN8l6L3k5Zh0LDgFSMDCoiGFW+KlVFE9xqfN41k4PTvbR/ep9vOBbxA
7Jw/8GWBnIsuWw2fX/GYOz1oHKNR8q8lB+kI/AnMlITBCltYkwbQzM0onLdYF5OJ
e2jaxwjjAkPRTzn6UucLDOqiQqzYEOo6jufGvEpt0jcy327DJDeOo+GAl6K57NVA
KkbsOin7ku5tr1MTAjeRxUbj++N3v8bGI2EKhNeU3X9Tmhq0D6XLUC0i33sHKswQ
vrIT02/2BOW4y0XMZYi5B6lgZ151wM79CE6/tUU7ErmntcDpZS3U57AiREkP8mF0
zgs5Q+komwXHz2KW1F/l3UbXO4hiVDHWvHQdMI9VyKSd4tDGr3trx4gTx3Qcgsw1
KIv45/0xAWceTBWVuGIjZnI4KxUC6Xx5fZfBJkgZ20b1q79cBLI4sNXFzJ/O5F4Q
50x/CPS7w6XX4uw+xkqEhXtYCTdO0yCZNSoZITy4762JS+jyzHi2ter2fOVhho+G
GWyvhJKIL5EIj6vQ0jWsUtY5aTqeMxMCbDEZQWB/JnXdrPvtOCc0lgTtZiKcxBf5
Csd6uNEtXlOl8GfM76+ItqDwZv2P94mKB0NrKw+bDkszjbKK02aBXyplVu4Cz4LD
BP2KJNMTI0hyzXubFTpXhdIcTA/bX4IwV47ej4hlFdULTpGh3qUIAVY8opd/sxGs
4Aj6Rz1bsXysCxywpHqy3fBSuC4I6TS5jU3O2/bSRJWZYPFhJx9dxbyvBfUjApRG
tNi5rFpOoS9HUcMuogXMBnVzSDNk4j3QAfzYq9uSP1nEPtuMwH8yl/2isfVnYJZ0
3iViNe1xX3G5amPsu7xZk+CqufHAQAGO+/iO8DZgzYMLq3GMhF8HiaHb1OIwMSNQ
JjgQ4gwFzlYbfcl73JR65g3WFmE4cfk9iAWAQqKQRIxqFoT5Ml0Da7WnZe7SRui5
ws4OcxvVn1jjX9FRgIP+rgk2o6IlO8xk0Huppdf8BQbN1+Vt+O9EgeMps2Yxw0Lw
nsIK2SXsOxDcwsvCL553CgRPFHjGk/UgD8JizE2dRbrEeLT+rLg4WMYS1LABNE1d
zp90ObXPxsyylsezjv6LMPu0R3/YEh/C/Rnauk+QU0ZzzQRn/TKwcgzBjL23nvli
57jUuP1AghgfGimFaqoic+JHY1yey4mM+KAY6f6aJkEEMY9/jNJUCOTnqyEwb9qN
2NnARVf1pJ10ZonHHWw3F9dKD+JNagBhhQmszILQkFzSdg+9wBlYH7U0qA9xe1R4
TldQem2yAPrZpWWq9hQdhVHEODE4iEL+a6jTTIzlvNxh0Oa7ifbUPcMMMz/nrFkP
qWcK8a02GQ5pojbYWFfUdoYVxYSFJ2YLlGtjQGYtiAJ74OD9uLiatGxbaQzaT9l6
/U8WS+9bjRCPJ0lubBEqd6+3416BsUjIoJMr7l0ZZfx/Zx7qGZXzzxYpOvEODm3a
AgIqJkID3Z3YFTlKlog9q0+cvm/OtYX7h+z1h65b9Mlem7b1tHNT6jBQZL2XzuIi
XT2VuI8NWW0cB0tG0HV/l+GoQKYWQZ432bkN8jJFRaHOcCapXmFh3rFG7fE5MGrR
m/pN6p1bCqNIxmKawREfgW2jB6SguLAtUDvJoZFrvQtYkVcAi+W7LnrIDB0eitIy
e5L6FOlTdaHwS1CYiOeR/dENxKs53Q12VhxAQD4GKCOiajUw0lGrxbPndFj0DKnx
Cb2mViv9QE3mW8mI4HoZtOTlEf09MUYGB/nf6M1dIi92bECm5LaXyB4CSd5uyWKb
Yus9ZkcrgoLEzCWlW4mFI+Qfiul13Sc56qcGNPzGFXR20lRzlQ8TzfY64YN7C+Qb
wFhMuTltwMX/TdBqWPshMRDJNGdyeqUHCVc6l+Di2EvU1AIeOzlHV/TfVbTxzqOM
HRgtIk0YUtOxJ1F92B2qwXwHrpxJetatR2c418GBUveexJ25VSHC1UqrM8occQot
cipvuBa4kwv6rTmguK8A9zuZpoye6EK4Ypl44gGvCrotU2jkJKG2eeenONp1AamW
DB+K3vmXl6lTBkecDHAm/QiX4YgXUAkvkruos2jFGYzvT5FxhoLfUW9I+Rzqeqo2
DNy0k/ARB78vDmntJ+u11dNz90nzAsg1Cr1KjksB21bPHtvS8QyybBWyVwawIWbl
ZFO35R3Y6yUjh7EOPJSC3JXSKiuCVMP0am9iat4C6nyY2O7ZxHTofet0LCSZaSs0
AklOYcZkfdHOkmmpqYARUoqLU+ichdk/eAmcEoY9umFu6rwxJSTeDgINX6qGlqa4
peF6pDCdFxPWPp7x7bTav8N3NK/QAovswHieauSfUkmv/nzcZME978vZn+uoZQzP
NyWmbGt/as5bew4ZShCYGg0OHrfzeyg1xIN43nhKOj5L2/nFiFW1yX4uX6ecvTBS
pMNiRoqSHjJvgRFovHKq0HQaCC8Oo026sUt7ViJwWDB7/VkJIk/Wn2n4TXbftW/8
JEa5deRRHUxeiNvpn+/Br9vXWykkbxeGV6TKFI87ySJ0+t+vgEDzxXU3UXhE2uEz
HqnDAeTsIwQ2HBVebhMGDhkWH8z4h1lZV2fmluwuY/TY2T+ZK0AZkxYSAeEIqmyQ
FYZdrmIC1Mo1hZabSTT/BtHYfA7995PzMHOtexewJ806hjML4E0RnrVzDx3uWFGE
AuQZeqw6QqsubrL1tFvJDYvbS9pJMGsZXop7Sc2pmJx/+AGOfbbR16RiBn+cEvVl
pH0LcgY3Cp/Mjqx4V83gIkzMXEe2XlwvaVfxABCMbhedErvm/WpcLdWEYnLeeM9C
L3qDjuqw9w2Ru+LtglNFszGz7pC/bPvcBQDbESs4P0b5xyVJA0rNanuuSjaF5v+X
flB+2U2xhrEYcEGQWpFY+MaJfhjsY8/MwkoW/jDEehvK4MVQfWz8qKbbguFJrTDk
ukWJO+JHuPaLaGXeaIqgIIsqDRXOhmFhztrBvPqkduAGe78LoI+uE8vkzMk16dl7
Ks/2Etf8BJ5+e9pKKD0UkJY5ajWuNgFkPP1fQ4QFsvqSH/DkPY4rnjqtvxkoJIrE
4znDJj/eaIMJ4GEj/xT+sfKIOUcMu+DZlmrzmz1W7206nwc/igbrensXpBDscr+S
H0LyRUZD4LWL9zfDre93S+DUcZKWTbWO/myilO9YGjP7Jz6zQp5MX5sqXF1mzgLB
9Zz+0dsyiXMIhCuVsrcFXMeeD4hebYzoOB1HErtlJKj2nNX9QrIUFQrlF1uUYrJZ
oNyDH27NkLrgJ5CboEAw+coWCFzIKHmS5yJB6lcA0/GxiDhciVcDGrSTEbJjCnBw
N3pWlxT99lRS+zYEsf+kW+JSqbnMYY3zvjZg3XNRIsqNN16C9Z/cHnUw99GriKdF
aLHW3TqUhNu5UscqSXIWoVfMG7nqjFCMtPkqpPB/J+vGJIPzmxejMJFimybqupeV
tAVOXSSrQwYBiqMdxGP7ov2EzCar1/FyuOm11u+NkLiLaLoP3wZPK20DYZTQUSNj
lF0ZRyjveaPbzugV5lJNrYxUzah6UQNumeS1LEBwGo3AMXLBnD7NmHarvJ+r3GzC
F/wArmWEB49eYuFVWG0v0g8wi4J8mflSo0aiZ986LJvgYgypAeK+7YJaPS4h5CsA
yEQ5N5pVoFb7Sbige6p8GDrVgtIoK8LUuqwXwRXm8WHg16fZtmNTHanfEYrWN4p+
MLli4q9SAufupij099pd+4C5I/DebdvVGpXbEr8uPcacJ6OdswmKu24qDJy1KGj9
F2L4bniMIKEs6pAYkBZxjtORCuysR2n0BfZgM4A8EUCPNwZC7pwew2RsrG0Z/iZf
BqbgziIPkx8LGecx6yNc+SynNlzytKnf2kCX1UeXaRF+h0oIgDXmXKTgsty8y/S0
3Q5QpAmzMp1jn5HrDska4x858//yLN1VDvc5DTM7R4ELdFQrPgQ3XxZOBn3KW7pR
9L54cObJFS5PvzI0xwgUwUVH8vJDRGnM6PslKSOPWM54V9hIlGbQVwKKYAE5bjk1
OjY64tvcEElDbVi7Xxya3m1A9vixBZKETfB5AHm/FQX5xhDV5Mdo1khesO6HLGqQ
U+yoPFFp8hHc57giGj7roLR+W9XIEHOmDq5oiW3tGu9xNCT9NswmU7wTnt1f+T1J
hM/0Snv3O0UOqP7ISb2QPGuwhhkEq5yEciUYj8T/R51uDpgXvZGYhIhksuJNxs0z
5SyGccsaY9EMkrh1FLR6ePZLVa0d+zegIay4osfvYTJAbFBvm56MxeW7nmcnEoF3
VsbjNaggwNOKhLxuyluVDIh1VH22sTTVYnTN7G3dANnx1IkQFohyf0geb5nK1MXm
JVJ1/zMVBJ5hfMqKFWp0a0XMG7c9DJMNywKcbMMSCTsXILNp7ABvwD0lfLDU4qJj
DCXxbgOjGprHE0hHGRt9mKQUhfwtvq3Y4tDUR668DHSw5FNuPnB86/dXo1Vgj8SN
SujDYCS2CYOtLubYICuKR5il4t6BY9ibfUzjK9kIl3V6fJIuDEpTKoUKkC4O/+Ys
UYcYff2tsgSwTskx7GOyJCQsfTjBNlAvFY0dblm/lcDtKIefj3ZZKmPEQ0Vwjdy8
s05S4lXKLORz/NKx7H3dlU6ilZmyAvJ0sfJGnY5wUBq8oee+oPwrfZw2+Ty9OjW7
FvRoCSyelSnHd0mWr0WfdbkZkyfFzN7xwW5cgohP/hNp7HJ5EgARb3hbKXANZ+6m
1VRmPyvefqN+090B6p/hOE6f3L8/fetgg7nuVuR0SJwswL1Z85XUqbQldlZmRRvk
Bxfd0OFCweXGURIkZ0Migi6fpLBFRz71yBy+Yzuk2UxveClYpuPYKg3kVGPBnZrQ
Y/MK4mBhsNCGMW0Kl4x4yd9JpAGfRrdwNtGtKu+XBi+DLeCUDcU6XPVm4lhzIsNN
z+nYkWTPnYiO0afUt6+zQmFopOirvg2/WnCkUBWEqzoHh2281clAE5fmZtMRA3J0
khQ8CJC/qz+2/Mx8OrL8028EhtUcN5BQ30ltxbVAn8vCL0hiNuFliPdiAzFsyTc8
ryF1Lfr7i0H8ealb8af74q943GpTgDbiMsrtu1itP+1IIaH1cGioTScn84LHuY+c
5xXzifVZtJIWshDIAtMvUuqXd7LtUS1Q4hPmzYbZmawbk/U2Ryl+hsm5fIQxa8wp
NhBTKhh0HdGO0l54DUwP1rjDKDLgZKdCglx7QCl22lhFhkgKFL1y8tcnAHLLyv58
w0gMamzGM4HGxHIJspyizAQukHZE7WSLaEb4CyMWm5th0LmY27e9L7/WYXqUja1z
/Z2WjZm0aHDY18rGP+7cv2nhkRm868z0meRPe0v3Xm2AGayTyQrt3/qdqKOkqdkJ
gx55GDtx6RDp7BZUE5zi2fH+xb0K4ip12NzYxC1y7984tnCNMnF609bMCwoQCXN5
fwrq9BoXwoPg4ifen5jlAk6yI8F0AURw9nFwzzzQPgtg7v725No9UQf8iydu/d9B
5ZVif0Aaqd6h4fnPZr/h+EvRHPPjcbdua1lHIH548qkFV+xMOCFjkCqVyEhOYpGV
sNDPNE1wQqJpkmrMxJM2JIW1L/Je15VcJSVQ3yuAR/EDpQyvILhaOZEJVIeTfyYk
kARVBwsScV24Bd0IBWMTIugHxPhvzrXreiHOgvHZZpCcC5SwnIXGynWEikhVYKRW
mVuGXjli9BSoCD65YURdcyK/OZnETdi25UUNn0QvjGPk6x4I0fkKj4NQwvdeKTKc
3kWdxCtFAaKcCl4KICuHQXXppB3x726kS5ZVRXErJCf28+wxXWBIzI3LzNf/2oDS
fYu/ZMD6jVua528MSiEg6xlGmXO+X+oKIEG/kWVEEIVT4EqDS2UpXUjy2btZxbUI
1OxEQgzWldDghVwaYxE5I0q++kMIwzQ7k9S9l717XbVMNxA34a0O5d9c2ATlUUeu
qJ47F5d8ykcv2Zel/GmrnTMjL6JuxsNKEFZ0PmZ/jMz6wA4gJYESq/DPSQPqj/wf
GUTOTk7f4JN4nQ+8x4irxV19oglyozSBrCe4mzIjiHyUhhNGXbzJ3vD1DzPR9i76
rU9q/GZe0RJt2aGPw4FVxosT+vj9Hpl33HpBjIvJ5YHPb7fJg8xVODRfSvYFNfQA
wDyYgiY/1f7XN+Yjdr4We5yCd3XiU0YCBQEH7ZMFXq8QeOnbTdJ4vLfSK6pY/fHu
TfcD1t1prt8ueFIoEdcq84hborcki4593z4lkKjRZfyp6IOcWCSfw6fJH+7TJrpF
yAM4KcisY8bK/5Y+GMfwQ+OFn1vqpHcp9EVjS/MwLh7L9Wc3D6f9OaLgoj2YpaOm
J7FTh5W8+cucCox3mwLJ64LP56TPlFq3x7SE3vh9tWX4h4CQ7EksbxvhmWE0aRWq
R6xJ4pMRYHgtVBJBTrST3G94krJYfm5Ah5/xTp++v+4gsSlgESBYzfWmAHHh9Q9E
sCtY5dIVxA4uT53YNuTEmMEvH+3I5+k1WhYHJJgTH/ZI9qB+xBPx85cyT3xExwK5
V+X+ZBa+TykAR/CRrrgH5omFoG+3xofwr6NW0588y5X22pQWYSZFsz9VJCW/F0Bg
UhMVQHBZjEpZBwzJOhfPWMx6t2N+F28/dLWOtTP0GJ0OMMytvDwYkcR4n48SpuST
vHGbsEOyNAzBMbfZwjwhl1fFavuQGy47K6DVwShPSvhcGX0cn+F8wOqWP0079DNy
YmkZldfhLgYiQpopJf6wV3+CjNvk5rywRLFNvWBMrFCdTBmDc/awjb/QtoDpq+XL
4ioyvRJUId9XlRE91yyc0DsgRjW9rdJKrY4JUhQU+7es1xfRwd/EBcwSqfhuZDAx
34UOiJ7NLgfZTa3OlwF0OfKb35HTyHzqovFtcT4vqct/s2Am91lyWIaelO5wZn7b
G9SnLM0Hir6LeDqbhz8sQFkW2mUQTEUBO1TySzcNzrO/1kyJQIeHXgiXLVM2MW09
rquQynRv4BaOXjLZaKmav6x/FbyFqBcpZgMhH3EDL5xOYG47pson9hAeanA4KN9F
ZMYt5rY8r/bBg+prmMXm08FB8RI/ap63rYkzPTLCCDXsetu0K/5ThIobT0nv3PxC
ojv6ofQ0eRsajmK6KhVizBiDZFOGJdOsoDJyguOrmSLLRgu0EGzEvatNc8h0kmq9
A7pIzZBcCKe709pIXBXlnHNu4cn0VCKCIkt3jxcKWZ4aYup14/49Su13lYSn+Bft
rrsgl3eOLBGvBNy4I65QqH2tGkhcDVBX26DOd0+99VBaHfxdbj19APYv8u3AxtGy
ZSiG+024viuFYcXxrqpHdnyx0vK5QPmTGfkV3Kasq4nPqU5bVLG6DuGY2K6kilY4
MQeH/KpRyGbSDRdBfHTl+E3gRGSNHGPJ5S146Qed9DISHpPXPriKEYf1b4wHSArE
RE1unOnabyFRmUC2XbzZD6sle03QSjgkr1YUgZK+5XPiUDmt4LLpDc8T3Ux9gCm3
T9xfCCI9UPXgNuG2LXHbRddGKRoKeZEr/7CxJG2xrQT0cjOrsD/NC2l7JNhZ9Seg
7JSl3EqTf8tHeaHVVkGkVBsYGu8j9584RAWc8X8AKn/Pe/oqcWFeDm2x4quPa+HS
f8uzJhPiNCIUN+3Wv8xcVPiHHKql6iQbbRy2qOdCLji4NuAenjRCJYu/vT1hPrtZ
BX+8LvwqIvnVnveCGzhzZcvppBaUzs7XgydKEi0jwkFOtuSXl0v66wOiiI2OkPoj
rVgJV4My7mISd6QLt0PCsajkTrMHmsZoETOeXA3hTil2YVBHeQHI3/AHKpvg76Px
N6807ZQEbZNxFI0tPf/CboglYBtW+ciy6cJRJ1GA5Iltm9dlNsSHMxYe64PLlM5j
ILUKtdWwRN7uBnV7kj1vj5SPdmTxb2R8e68cM+sH6jA0mBq4zl5DfIxEZBa3A15T
SQWRurCNXrneJEHMndrFfcfwLfslb4k3FNvchklxp5X/u+A0/9G5uLLC47KoVI5k
mKpy9EfhZ4pdlGs4nnsMkhmU310NcX7AlsEfbx+bDhBE87yPa6XQ6CMn68bsyeR1
jDwuY9gwQ4Ss5yiwDGGEN63kVFR/x3ZzXzCxrP/zlKwQNbMFDXTZqCzZ/AfknU5y
fvvCkShic8IgHEkypOEZsWMT41uno9R3Xkj6GPI8U+8YFcljTfkS5xjUH4PEUNEx
YTrzeTunCdvjqCbpzL7AUSBjlB4Su5M96uqHnncjBC7uq9a/MfnzZIrSPXS771Oh
Uff6+3/p7lFzdBUNa8YXmfIfRLvcsNollOzWxmSpLwIDezWFLqtlECuzX8n/QHdn
luQnaF/tSB2ms99hsvnPrkmW1zd+m+WWwG6WN40w4I+kOY323Jai10FWSuBzMQmU
UBZ4fFyQoFybHMC3/+6FxhWx/B4+RHtRxx2cPD5uqwhWA/zS3TrfpZc1Wthc2ecY
Y9zeKaOrh2ht69PLTF56zdL9/FerMdjtfbv98TWOCCXGunhcz44v7dcaB4w91M9p
J87diJ4MhpdPy4H2o/GczJ2HgQwlPYk0PVjuncwBESKDCtR5Fo8/4hHMgx2cd1Y9
UW/8cej8eBPveeK6hDE4fxENVEAPiURf64IRuRyY8pJBR6hFKit5Ojl/r4e7bGqX
5JIGM6itLg0rmkQIjMI+tXJLkR2B6ooJTy2Vrh24DZACNFmYHE+b+JXG8nYSXm9n
VTdF/KDv2DF36SGu9BKZBvDU4e63ZSCUXzbzx+YVSnAfi4ZrbrwDOxTKT4kyx0bb
0e0eWdlnRumPLUZ851NbGJAWnlort+ZfBFOrv/IJDwzWoPlIgRA/uUrZT2k7ZtoK
kZcsq7yi2FFESDDBOjNUfW73AqfO/bW9eJBG7CJ5TTQq1/vTwFWjKjZk619kssRt
22zFwyilyA4tCDl9L3FeduVMS9TXSOgjiww/JarcxYwa/fRK1YE9g1+druQpWJlC
NuQcM75TxbLHfjc7gcZ4oK9CShZrtl/tHAORUA5oz1VcYVBTaYyEUflbjlqqD/Tf
JOPkELQ+Af/tm9HjIIK4TniwpbxTr8EpxaIqCNoz/c7x7IIXQXGLE65FaWOX6v9p
bx/QucpA5+qlienmQZ7ebLXzaLPx1wgF4G3uHzA5+st3QM4FAszySwiuiZeXd4x6
Ih43Ney6SSsW99NfPph4Ne1lskfsevPahKyRxwa8UXui9LMeIfFQbXkvv+3A3Bxd
CPsTreQ1aduKQC19s9FZFWGkp4sPN4FZC9Tszuc17z9cMx93xkxSAl5gLsAalQ0s
9GW/8h30YDNrn7C0X8CREg0eQMy0NP3BLsINVI/UoQOthHCqyImE4ao/upgaLJ/d
ecOR3O6USfHypk4GoNxB9ms4Vp/2CxvRa2PaAvzx6ql/17NCXxbasdNkErcZ3TAU
sip5Bb2IA0RIiON+uUSiAeWvND/IN/S3tAQiJ/qgiEGpcXgbM3aLeiAPS7nBkvPX
NDcDiO7f61dPnK4QuESweypH4sTm9DCfxZKXPRzqmEyXvpoidZRb8YkAqhtQFx56
pBfk2gOgoDp3lLlBmG21GjohvixckbcYSKcGkC/MwWVYO9JT2eOcYT+xd04f3LiL
GifeME+AaiHEn41oKR0jrOZQ+tBeXzf7cz3n1OlzUfrfNumoIga6yuwNvqqQyiYr
M57qtkP799/ouqinvh4ByJcyrrrnTfVi4oWv7GaTl3ptrccAIFV9rqQ4k/FtkyaG
k/qaur3WWpKgEzcbDoWlad7r+TSewKmAwpyycpn5K2OM/DDvmBp0HF0nxwsHgFoI
XtWIOs3b5JnZsel5kIwTIHyBJ84iANA9gXSQrP0/uBgFrRD0h638dtKVwy8j6Wc8
IaKUEzSIY3En7swxM9Ogu+cFvFQAte1SQojYnUFlzamewazw3lAySHpHMFUvoQ5t
hiCa697GSstPWWje0sQoxJGwxgI7YKTGFIeuyOKqRZYFdamrR3OmDk6jDCRJwA/i
zX5fExmHhzU1eQRgyvhIgOVC7uDy+KTNLKOaNGs7CWDegKWWQcxsT5evVrTwcnLC
Fk1fzYW+4FzqSXaM7WmV8fLwXAfS/xVXgH7zIUpbBj4Bb0Ob0B/JJoUp1GCwTNbs
3F/YXUhZRgTKfoLFJr6YrBVYpMUwoyhmwcdSa9a5sxkavnWi3lTObyi5bk1MdPBH
EqqNHsdZVU63oqeRjdBYRSvvzw0NM/FPwNTiwPUFkE7dgdQ3AkljhSq9Nh04khmN
WaIyg22H0TGR7UEeiSwRtBjR7sC3tNn/eoVFLNNv4G7p2w1tRg7TeeL2zLJMFF4x
z2Y879UsmxF4RsVU3dGRohjfGUhqLb7AJBYauO8d0IIGZbgVq1pPQETMOX+8D4+9
nGM6rN2ONerQ8+8p+REUJh+cZERaIQZscAJoeEIqeOooLS4Kjt7YqfguTNe+SnbJ
9FrKeWl5CsIYJj/RNZ6jSa8CtuQU9Pe+JiVJj/nnez4bewIEhLesyI6Y8Ihem2Qy
8uUt/LWlXWvFIVm9+Ygf3RKaywBWespV+P7t0LWjfaGbMbkBalT3OigJMpBGaxJw
mhHyHdIeZRxkzxlwgs6Pk2DsSmW8P+yf0vY31/0IHsAfiUp/JzJX4C5g+H+5hoZq
99SoiC9t7j2lrFPUIVWXeE6mN2R86sGZhBrj6hFNN7tVwD+4l2w7dLqqhVTdf5ml
3+jQHRSbIDZij0VivODMNTaOPQiTiryQDXJN9s7g+sYItQktjIr4vq6Fuuxih8YG
SzngHSU2cw9k8NmKLnXWGrzKC1M2dU6h7WMYQ2Rn/Zy5f7y4LBwrYOEzHEcceERj
YhOOF7i7Pd/PsxPwe0Oq+GTqoJcaWsut3X30k7TvOY58MQtgl98BIFmGKasYr0Pe
f8do6NQdzMYNcqv8r7cTGVTGlnCGMoKO1bqGUzpWL/zgla+rSyrXVa++tJKAP3VH
5MgBiqaI4g6j/W8sKPAMkZyka+d5wLmKdLyPh89FRZeZ+/OgRBGmH//IYutGevlB
spCaMzkm9YicvncJlJ40wyGJLhpzpKXyiNXz6iOblAINuMS5EM3LP9US5IQOOZUF
nJmXSOztwmoQZjp6feEsh5cw7XX/j/LNuQiNCADNMNlqJP2M5laT+PcXGnPMgI02
VxcgtUwWdnTyRKIsVS4CGs929dLsLAGhjJVjaqXIthxWMlBNG7uN0ZNMzvnP6YeT
7YSVieP0bd/3LTI2I6CnAql/BYZm49A0W1aWucQOO5yTIJNJIjK2ZNmOHfXa8p/a
RlXV7FIho+l+W2c+KfCFSydRGTURcpFQnLdKZbC00kEtLyBNGDw2eON6XDAfqcQz
PLWgC1bUUQD+iMJtP4O9Oe1HoobYafp4ND2pJTaymbPVSG1JNfa8fdIvd2jPw1Ni
Sftb+OEODEeuaAKPILqrEGBAi0OZp9jFfaZX3rFjU6Kl5DURbRhPAuIdTVtjJdsU
If3DI1hlEVUIxZRb5gVbIa/IT8aszRjyxdZUxp4Tf43HkXxYIqV/zKH5kIxuYmNY
0ivXuV6wBILfcJD8Youlv9amJ78yCG5ICv+xKGdhW5ZIFwdAAPysmq864M1Z4z8G
g8gzfIikN6yjKQNQzrcWWOITeLlSL0XBRlWBvoDZ5L/vUdFpt5FcDtGadQPONnva
ssCwkl5+p8WxLSAZ9i0yUNr1+gOI++DWT//YsMgWrjqxIa/33xY8pv9OtlAMJ2rx
vUpyb9XiQ3JOJIyuqoPE4hgNv98vYI6PRXMgS/CazVJX3P6sdvZmnoJAkiZ4wGwT
SbuDvUaPuXS64dUgG+l49nRu/CINbVV+G+X+pd701vQw0dMRPSbTnhbr4yvCU7Vd
kx5e6Jj2U6KRaTq9q1kI+h+djjctGkVUFNOSh2n7zIKjA2zS6LTRaWLVDO09BIrB
VL6AdXYFUIklGDde6H9/pA0nyvS5lQiyp+zBTqzQ+SvKanFePUe9qtdtW1RDu5q5
vtQX0iW9Hy0+qUN47Fwc9w21bPjOpHHAOsJwLwwQEEtrZYAVl6TDrERc0FtaPEQB
RXnq1iMmXp8MGQYlcm5ibAiwnWKD+3rnHiDwlGNkxAsHlGXNLenOnQE0AKeyRUb2
rXUejjLphWvr3vuOM9jw8fLrkylvouVwlICcKcp9RCHCxhIw7PQKSJdwyfq27pBL
P9hVU6t27ttkRvFyJxQWB7dlgmWz2bKb6bxlmK9D7gKoHdJyzkWdt3dkPRxICN3A
8LDvWCEoTOmeP1+MjAoQuG6EHwgApWakvURAqnKYPmuI00RDyYSZxk0r1z57bvR7
S0atkGM1VetDJiXhN24WK6ZGrsTf6pjDK29a7xY+J83gymYoU57O1CxuNLbK9uUU
IAW88p3yXl2OyxovXtDQNuBhyrR1seWS8lGgQPWPLekwA2l5W/3UUS60oglMJqe0
TPKre7ypFDdqKytvLtYk+T77ImPAMO3sdqpwFuly/SdoNJW7+mAPzDoWuZ30aFPr
u5N6Mzn0rduKQcPvI+J5Z40N0ntvxOIShiJNCht9AWvLMER4DQWvbo71ZS2Ebejn
+lFGHBm3X6SaAyFKvyToBWnCHQN19m+YO4I48ERduWpuVFDE895VnL2YSzfape79
Z57THxhZU8aDopGgOjfMaD5NrF47Onnrr9T0/Nf3EAkhe9D2x0rC677KT8WRo2NI
yPDdcq8dsn04PM5HrM8/u/PLanQ9VgvMUIBn0b02PVKFtx9aSrND7PLVjqn+f33g
wwxJbPUJrhCfrTOyY0XkKDYFqR350PX6scD381fhHyqpP2Pf4G9eX04EZKqtfNok
bQdreZKdk13xnJlEZ/lSqD46PIbld5cibsigyvdMiZLbQ3Xx6ses3uD7+XwSQQV+
GqYorVSc9qAr2SswidqVKyk1qHuCMsDwJgUtVjFE4rDMRmXGcJ2jhS/eIzTYZtoi
nzE4edXYi6LW4SaFfIb9PMo8+1CdSv6V9EgeXurB/wxApf2gqy3owQbDriuH5y9g
OPnu7FGwDHlKRRj0yizRkcKZNfAPwTiN/RoxSRqwq9bh8QpZfC5qeUJXV92Dulxu
SxgVWjzR0Izh+Q/vYZQDFSFkaY421S/sJtrUVF5C0R/0GUxm38nhM6eLoRnIB4Hw
8zCl8ksdcAtYLGERuIQCCT6Zlkhc8rkfoBLasoBaarSQu+0hCSNJ1NWITg77MTYz
K20qQeG20zrBSq2K0zpPBj/PET5DTnw7VnTQRb7vTEypdhVnBgaIRSer8E1sJZAx
vVtMjPOqmNyWwky/Vi+LWqLfjirxQbhTgq4402ynIWXsJDOPBeIyAWc0JxUYflxD
1l0XTLXpfH4ocCXcoAqTXaQcfj60KFFmwkMQEEquxW7v/xmB84n73l8YlcZztmnd
5c25oFGXqd9ZTciGf07WM1gOs5VhKq2hHFX8LhcPNh4mVFXsBFYfK9MsT77IVaAm
qgsonekxNm+ewVqgwMwEDCfh3kM7dYJrSWQTZTgYOQRNnTD0Etq3/vadfCb85M3l
s2STls+lAWADaOSyLLrikFOHD9DiLkdQLoLGIJ7D+5BWEB7K/5oKMDvmnFkyWZuy
ejMs6CmTTKbCSYdBzIkUM0Vd6uZ0jbcIWd4U28U1Xx+knYPC4Xbld27DyQn9Jyks
Wij9JWDX4q1lpIecU4zjwQtQaH1zxB1kXXLfI4JTcF/LXPQGHwaaprK2wkwRgYD7
BrJgXXuhYaWVDLFUbuAxw6T5FBe4gDGUM/kYd6NPz+LhB0VF/8Q+TNn/qtqXiQZT
HKr7axYZapN/hSY/S4wczYanyubZ6bEdnrBH2TDh5G1K4Ez/ozRtQuTWVOiC1I+e
6KB8uDqqM3Tmsw7QscRcXQha/rDa1UUz5njD+f7gnyaelaNJY6Ez3Lg39+FMUbTe
I5TyNxKcPEr2Id/hDd+xbxfU2F9xiHSJjJYzrxPgYw9jzvqU0jgT/9Dvy5ivLwy5
MjPvC+uxAgfjxTDgtokz4VlqK5yoqs8JUOGA5AosgA+L8RGNKmGYFJ8VFOEGUwgU
+o/mZgnerStmSe+hZYpMTYsswWHrFo+5Y0e7p2Lh8sXx0l+VOGNdCiBJmZH6uKmu
NKzZPpIOSJarrie2pCEAJ+DhycDr1B/omhDdzhZ45UACqa5JR3iK4wIlAromKPUg
YiWSAnsJUJkzidRvOAOAwHKKRAW5HoZEb7Ui0YiI4kQlX27Mtu7tGPeTScsfw+VX
m9VROoOaGiZX1VWJk6wHNEPTbAUL7AEorgR/WwXqJZ7j5s+d1/Ng2ulcmqS4VSYJ
nuqZTA9DdEgstinjVF+bAjDgoE6fN78ka/TXPAjSICzOSPis3fpDmjPvUxrKidl9
pgBeMZ7q+4M+SLkqptIrxjqcJLgp638aDE8BACeN+4U2LvGZyRerBdUAzBn7yX00
q+q5YskKdChdDxNYQKCOWU2i4MovpGz+Nw+khorw639K8IWJ/9ngVnB8NTBwtg9c
yuhsY2WKcQMs2Y9LFakgkNbHrojGI6bA0Yx5pn/YFiTWdvCd9iZ18W3l/+71eirg
sfC7WbrHyErmcLfh3BHvfS/0XoVDHxHer+qqn9F2WNu6LWXNnBU20KpD96oVAZmJ
3u07wSVeGLhxGJ2c6YtUT77qMKs5lYXfSwy/HqeAc0N8QPGgOc5kjW1c4TyUPBQw
XKMbIIjRvBCKQSvXo00AOccEe9JThyRdNA+O06pqZHcvX1NhGkzW9HWvAbmFglRL
T0pg5E3Ey5BBtHgUmjN7Z3YUwBHAvI6WbYmjtLavJNCNcuUoA01sGOMh1v7ZnzKr
P+MLQbaofVhvh8E8A0eJkEX847I9A1LIdcURJr6V/qnEaYnEXM8r2rWPllDWXfLF
Vg5dZ6Gz90FpIlIxOtJMp1PBvmC20xFphfRhtkQQQ7nSxIto9sOoR/KDc/3wcTYV
jWx1y5Q818YrTQ30hz6IAL3L+p27hlI7a1ZC4dve/CEkMMFsxPN/MK6zIYjHdffG
reEPCjy9b5nPJqTMjRdGC0UXvYQnIlW8QQvHJs8VF+fXtwwVYH5kun76fDZlDogu
Hl/xz4x5ndkMWvbgCeTvxdyWtL1+5It3m2p5RGetIV9NYUBdP2txQRndZ8BnzbZG
SuIuLmgnD7MStPoxQWc8I2w2Z+lOHhFCWrMzeI8VCWljTgtWRt14RcMRv1C8Q6Jr
mY+RWAyjP7tc6wKHAk7DbNe9QoiCkHSqDxf1aCtHl2s/8nMwNefbL3RA1g4Joy3Y
AiIpBVKLGuDtrz9aIgm2vsvDPQkgM3uHNkKZKRJoSniyagGQsaTXGLJz+obP2qlL
Zxz6dsa40bNLZkZg/Uu0zRk8Umyf6srJigMytvkDOA3pAEc+2ESfHv/boGVhSC0j
SLVxlO7FYBzUwfpxvyMfJJ+8gUks2aKzfTMESEORvuQUCrD69hPdEDOJOcHPfsr2
Ik2C77rJVK2ZFNnrtAsvig0of2mWvkQVRfwrs/5VITVemVZHhcEI8DGtKr7nPePy
2/ItP7JHaaIpaUoDDjXnuNVFB+eOuOChHJbvQgeMOfdqQOC/KfSYBO4+u8ajnagm
zyOHQHK3HI4X9baEhGbmDVPuvNJgI7wNYDIYKpEcZrAFaV+kWSN3yNO0BBXLZ/uj
z2ADIN8CiNWz/3bnmWxS4yBFf6or/BaF0INK5WYRgJ3RkOBCs+eMIhXHRGZHemaI
a0TqPBryJlIMom46cRDKzrkMeZu5I8QwXLDdgD+b6Wi9+PLwoMtFpo8drEvD5BLs
pIxS0+gN/ss43tjiZ4m+tLPhFzrZgZv8jauekCsLc08L0nHHInF6TnkDhUwITn6s
9NKScvUIJtlML1MYwTVZEFRsSsYWO6MYnbNjThSOAjRCFFJoK2+DwK/G32VR/y3O
y6yXbFbet8RVKY+vyFvj59sSk8sRBltOUM4slF7Q+ynStBb6/tQjgVMyyLoH4IqQ
8x/uAl1VQ7JAavQh1Kugz6yJGUzYgR6b3y7q3yK1Otn/ONWlSeEt78kH7M2ggzo6
ltJTQAJBTCiG6/QX2duJUfO+BJ7z0cE5KFH8JvLGdDiB8rATEL2vgQQTrBABryR8
SMcUD6CzGdrFJSy27OtUp5+kIC46araJy4yBFLyJSBbvrJHQe2YYHd06ioa8Nxte
lsIWpmZQJ9rVjaawbB51f37pcGI0tR9DbMgSm4hRnHhCj/mZJgHzmcNrvXCowAYS
56pZpDOJNBC50L1TxzF54lqfsRUKXfmLH2XER5lLkkwKBy8QrkLjG5sVnVmfR3W7
NLNvNNzC6UqMfIzvubWTsKWMN+Clp88qLaza3Zviv2l4ixFAsrgw52GINA5b5YNN
Wf05TUrjA3OzuejWrjbyClP+9IbyIaJaoKW1VCfZQilXsexPomKDjVgYGp30FPes
n+G9UiCu0Pe+tUCIb+NEIYx4QS8k0B/akEvwWGJwCVMGkeNTEGWXjAHAZaaCw506
7IYffAnhzxjPxhAJ+AqeOBS89X/k0UDJrv2SxyazIT/NCfcv42kgXQrm0NmN1L6/
PQbBS+d4/tEDtlhnLj5iAe0IJgr8ZQbgwfwaayndI8XPN1mhKO+NuSj9Sf5WtHbg
r05ULEebdBpe0aaLrc8cKSlYNnu8uNRhCncWDoDUajSdHW/tQzMDbc3AaCiqXt5D
evRN2KzkRxWaaioXh/qMBInsEfO6jmrDRfbHkaSCJIlqahe+h6VWMLzjNh6wG19n
S+pVjoYeuv4mm4xyBhh4RoQ2+TYcTNYgHH8X07EqWpWoh2zmOu9VoKtpPztXSX2+
Wk2ptEMpmTlLL1l3iKSXDIsfvwkpQrOLdKVN5sNCGxWxxe5LQv5GY3AVfSGqx2Ff
XzHnlIkRps7e9iC1ismFAJTC8lozhyo7j72up3B2KFinZ9GWteumcUB9egOSgOna
PipoOCqFOuN5EpaYJzU8HwQpCQ6ZgnX0z5igNWyr0DLdWXxM0zx1gRmKQPiN4tMB
BB5PDHVaogTiIiUqhghSVvjnD/fJev1YOC9/Izm0KvWFU56fR23LBL3SB7se3VV3
FX7VrpNb4tO3u2hfaLh+HYR7FM7ME0JM+gZQCGl1ANuAzvxqO9SDgIfEI42qSIlP
0aAMRkyXduc58Xvr+QXNxn2JGKPAnN4WPeyVs0SDgDx0N+dLkpDxP0dvM48BtJ7O
vqUzPYY2DJZ1Lpb8qDbVXK3xo8sH5aqIdsedq9umpR6h++QJwLghr7A4jU9uL7WB
JL6Uz3fKn04wMimz6w8LXrX36LO6eGclFkH+EfM5wKXybfFLhsodVs8ljQUS0AKC
9f1loKIaBIhFIeJatFp+d7ZX7Y7wMGk0F6PiXLP4FDIJJ1vMWU3idBngsGn1KDkG
kSvd6MnGGUy5/zjRl4eFV/nCplNKSvR+Wp4OmtvTTQF0sCpJNlNRj9IqWF6K/NIm
9io3fR0rJVU6AuJMkeCD1Y7+pob+mSdUZP57U6VgnHLptFWCzU+KZqCiAk5BJGss
BLCSz4/QD/RGDw0HlE6haGV8srzvFdABgqKmWQoTxsTeHtIpmkXaOisfe+BVgkog
XzcVIRLvJ7Y1N9pDmuRUwWBHNqpAb72kyP7gNmuDwyEb4EdhNcC9SUZguKFBICkp
Z8ccpbwGdXo4tcmYURplRyNPc2w34s/WsL8p5Ydk/RNsUYdFa/B4pmPCuZ7x5G9o
yCcz66OLtLUCt5VB3V1PVXMLnlYjiYIKt/E/xhTec8znBxLBoCYBsyj5//GOI+/6
Ll9DigFYi547vktgLfxwxH/N+Z6JK35xu1eAHqQ3hDbz+HwKi6ZwczyucuPEkX5y
1YGyD1lRSkRsALNdBswmNTShcEnfbi3jEtj0uQhYdR7x708/wURbYucKzJyvWdOF
vJ9cyqmRVIy/YE+tGd18eDiqRv/gYUn5Js7hEnIuw/RBrlUMABiwzERa/PQbxkE6
khe4/HYo9YrkqusJVgKlueKXeddOSX5HMVy78F+0LtP/G0uMo1/pVGlBzt7Zxyhq
rkvObdM5Cx8bH2TI/8WodE7HYVNhBGHgne9Y5xZne5zkfIL/vFv43+DMsBl78E1m
LuNVAIMm9ry/GCpmsJBWdwq31gOSUuSdi7gyeA+XmOA+w0JOiCYIymWruSHL71Ak
ki5fOvQd65dPepy727PINEJUIi8ahoYOeuCkz90sgTFXt/J23Xu7k7+g3Ieb9haM
WGATLIs97vF4xBuUzRkqmv/TIHXf4MhLmdoJEzTuluPks0NNdgZSHqQ2J5+Fz7gQ
0qH1s+Af61QGeL39ZCvKTaMG4tAaFFMhdDTxzzn5MDGf+i0F8HLTjF0kb26ttDxo
G2XfgfbVPuzNqfzEuppaFrgZR8ummAv0gdSYCoJHrNn247FzhaBzKN7JnIOQFqE1
jrkc8seTc3irROfBXBkMj938dYLhzgZAO5Um5tki7/QPrwjuibneqRh5iG6DcVO9
CpKkpj+9gm82UoA5luJ3BnBGc9pjAOtBTd1dF+CKvfmVshLEmEqEu6lXuM0hCR5F
8Q9dRBrz+K5yOn4OdrNPQ4kBi+QxHxU23zv5kvHRlCeA0fjzkc6eg+qxakXMseOV
cf+U+vW/aSXkBuKx1Gc1Wtbz6Or7BzYaWPOxH63lhQSFXpTiIrU2mtMOeMJEeiPN
dqO6x8BVH/nk6fWL0xliZfrJkieIT1obYEDc/M8qTyJ0prsfI3Ijmw8A6VW7H/3Z
hTsoEqGpBz6Jw4u9VHXFEJlSQyy5BlYmJ102dvae9oCIXBGm3fjO0WEPrAHUpU6f
s8+dxxdup1tTfgMNaXeh7Y04QjIF7+PQA63zCDktNDXcYo7ZSOMBoq5laaeUor4Y
BdGAiA3BwNCFk3tAavEcJTg29d477Gs07oso4ebrVpnxvlriFoEkvkb81HZ7shUN
IzPbbAuYnVY6XhaQDTLvgvtB9D+GPxN9BJuKHlnuZ+EyW3Wlo1mk6Ca8ho+AnHph
AmfaCslhAhZh6kW3Jyor06x3rbtLq1qa49Da8fu5a2VHxrsdSagnVK2fxBFKo1+2
CDdR736UFYqZyO4usavMCC14nPdO3gKnIdQypa2sOs1KjvXYWRErV7BwEOkGd6XP
5Acs2SksKqIyOCIDWzHnqiU0JwxyySGVUQShnHNKj6zPizCiVbnJo8Nmikq90ms1
K+VgTw1+jD4461n8n9uNoYMMFX+7J1zjbj6WdDsO/5VsJMwsmy2F1Nh424/OJUiH
u0K6cOu7arH9TB0IvbovSkaGuMJYhI/g4aKmz6A/RGH2SbaEuhoORox83cAtseBw
b32TiL2t37FMVJ0bTrdMRV+RpGJxL8bcdDCNZeBUbUcIgJxbZu4DkJuRIUB+5h5Y
kmcmenjrAAUzv9DuO7D5NebqlaYc3UGEvKtz/h3MF301I181aLwBkJkwFD/f2sAJ
6I/X6BEFNCZ5CnWp/hEeVa6UY3wxrgZWYF/XAk5yw/udeS60c6Y9AFY8IEEUmlTP
emlGunqwgwH+0Clls0zMdW/wrmDeodOn/DgRaGOlvUgs/9XMeQx7kLJAR3RTT0dN
A4GojXl6krTMfEqlm9uaINL1/QzccarwWHlFeHBDb1bYUiU/p8wwnanBrqB0vyTj
dVy1wEj1DDmxp2yCSLTwZh/p4afmcsNU2klAg+3PlbzovAipG+HSgaC0Yd8kLiaI
vgzVK65RhOjh3/viO2YICInCrKlsiKGTf6UioJTW9vk/VlocAUH9ZjV31/AyvQyZ
otx+W684TmK+4ZeUGYnqn7hKN6G0n4hetJTQonTIzXWmhc8kHxCyupRcVVddj6dm
RbOByVnI9z6uPl+3eHxiaZnkt9VUaixACyqFVu6r1yfid+5I/ra3NFUAOfmEErZz
LYxzxEIcN9hPOn9OfjULL6yh+izmHGDJE4ScjahYl6ggZS++4K5t3MH1o1bC+y23
mQJwpMTub9MGmbHw9bqjxVt5j2oHwAU9QLDRlqwyi+CceMB/fTc6Ywe3WeSt0A8G
6zrA3MnU8jWM8Tb7OAqQmH5rY4k4GXPkzqwDfmPXVvNnbig1M4ZqFNvUXJjdCDAE
lAWG9w89L5JFhDf3zoDnQ3VIC6NWDT9uyxUzRmu5NM2OJqf13yffARk/xN7WpfNL
c4DWBImR5kxgSi4YVu/mW2EOWusPLMfc7jyUpnSuVW8rzcm+wk98Cmis9EZQ9Cgj
xW1kSq6Zqp1xlak7/G5ezcZJu8jw3Q02ZPA5TRZe9PphkJiD29GogjmZnbd68yaB
QA1OnfAxiLcctKnxAre5MYdoOAmBhLoRiHQ88ubVkUq7gRMjlNt2CIgLqquHFlDM
Mvq1a/65LCefBfnSYVmYGfj2oYgYaNSGvDMRC5/YLxE47rdbyEfCWstLH51cYlTo
JTeLCTGnorWpKh7D5srgpt1rRkpHN4srSPmSMcGaS2tQw2fPclQ+fvAD+TMzIQhG
WjTfIqp8zqdBliAigU0758GfLRaQkWxUMaYAyOScwlgGsvMHHPoF2Ndh4wLjU/tY
A/G3HxJAYeCF4IMGC7ijj7wkOC+pocYevFNtosHcljEokT8ZaXSbo0k0mQmyxiLO
JK00HexGYXybaxXYAOUYRfvzb253Hfx/U68+nmct54zs7G2m1cBpxl7QGRC0OY/3
IYuSLtZoJrLGmyPwqNKyleu2mArZd6p9cCOwKau1+O1qI6a6lmFL9UCa1BLwOE0b
NNTTQaz5U7SAmpLO3OKc5sE4d18/1Bz/KMkaIvzHWrVLBV62k1+59UOxP/CW+oKE
1VOZP9V66e2NhhTRqu7Gehdhu54khFY+k6J/dSqrhWLeCmBtaDtxVcauCl259lMs
Q5OXbxOuDS+ZWJvx7vWnf2PHcUTre46kClrhj9al+tYrqbOaQSX/w0CtDID/T01t
Ini5yluvL7ErFz8L20bbpwOt1ZpXfbUmih9rVTcc0bn59o457wtoXgqZ8wtY5jl2
s9CoYQCIXi+lmMkGW1wC0DQ2zkI70CYUniXF/sZflkeDi9dhKtLPUR0r/Wnc2jpu
oFWx9blmCATkSCzi1IwiTD5vdwFpN5MnNuRuKwDrt7mvzmdbZWExZR7vxNAqL8ps
Yg7a/p7y+vl1UAyTWnhmasM2nwA1chZ0qPR6/BCmnq+vffVwMfS6gF/454xqGwu+
1UUzuULMGu7na5KYXtc7OIFbONTNd+UlAiXNKtODk4hu8NumB/WSKa9K1U4VFWC9
2TR27w+77WtiNzGk8F7ebiBgTExXoztNhYxobeVn/g8RRhHpP0D/ijkPf1ELAKuQ
WQG+L2z0U+myoghfS3AAGMe3z3uGOV4gBWyqmux6TUu4GGhvt3SYHiClhMtklxEQ
rHtq+7v3wPMTdbft1Ge9aTbmphwu9GLnT6/wMIMArpWmjLQStOyo1efeVJpdpjsu
X6AvU2WTZoTeTVyHb6eGGXUTQl3b9mA/lZYe9cN8Tj31FqHjK6fYZMiuyDyZ15kn
rFZ1+NJvQ8duOzipK1J3q4tNT7XxTTbsfkhcWPOuw9LuIM5qymQGc+sxkIx5qp0B
wbC8LWEvvaUBgddMAOL8wx4HoUBx9PHauY2A09pB1G0Bdmy4HCodQXBNWdMS+V48
/dyss77yuVkiELGOw4eFYnCsdgzVXs3B+RWrQX68YcjD4Nv4o4TfrshSvYAg0MSj
gyqGP0RdBsmSeqsI6oflE+zaER7buht2uKU0OxCDV613nqGKtVbiMlCxXrm+c/rA
NdbLk9GRRiw+2fqGXtetSF46imV+kP+48FKS9+ZA/uC5qubUFTr0iZNf8CRetuPE
zIWFfLXVPV0WW+1nji8jAddkjqKDNlQenrOhRnGU1FqtVt4G772IOOVZHN4lJ06d
uaQif+UR5Ty+rpOMk27um0KT7btSiscYoReXHn7PBpPa0h2ekiEN5l+4da3XwGTD
ioBJFQxJZ+wKuSwtkK7sjB2O3kyYg+eW5UmVbHh88nS6aSvLta8bLgkjARxm/f/v
l9/RSizfNe20RWxTNaMlZXo+la2kwwijC/DsvDOpIF7LyeEQZuxbnlNBIMyhCn++
G8DxxolhTh6okI1Pgtvo8p5Eh8O5qwbgwcWKZ2Hhs9WodJoUYSAghfF3oITII6QK
QK/Wk7nVtt2t+oN60ZoNgx7L6zYjAbxWW+Q2nDW2y1PQlq0748N7GtEh0AKuwcGd
sIgcuXd3jEYoRmkJmD63ODXvgzTVJDLmDHs2yA+bEutoRNNEO7esquLlyCB4BYwZ
DuuXmd3MB+w/bRWH3NttXaruxfNaP/ZOqTPi4sss5G1l4oAJOvpVQ0954gcAHAPO
uuGFkgqUn+EPnw8G30Bah0A8+6B4Xbl3ZPlG4WIB7EJ46RgA75iz130FFR/MuFfR
dDfcFOKtB1qG0Ueo2oWKeKfBxvrXRRYXLlBs1C9PQwC40Vna9EvOvI4M7+9pOViY
P6M7Fi+uIx5ZMea8JcnxV3nlFHzsUsFJs2V4N1T84kNOhbfcTEYSKQZm3TTTK/aS
VpA5isrQGzLv3Ht5TupQGshuT3ep4YYSUCfuZAQwZOy28nmX9sFOzutCOU9Nq99k
xnqLooEQNHorZq0jTDXj4Gez3OT4ycNS4B33PceDHY4IJp72dNvRd+lw8fdig6NA
eicKOCDGHSpFJNv0X0NL0kEkHBra3VH/5uDKjeSXI0UsIlRsmLnGiryvtGP1EXDF
LTpJFdYq3DcjCBh8eZocGMaFTEIQLChHXuYppgeySl2BzUXaO5e3pemg2okTQh1E
Z5NgsC/oIAv3RxJ9hINZeJ+qatjhBu7d0OShmKbg1h4kK+Z2JfA8vwtOd/pPsFP1
gMFCS3NEsHx7aQ5hjGknMBTn8JGx70lzPjmsKlTxYjhZI00hkiBRN3WVKqoF8MRu
/Eizur/IEcEy8tCOvukxtg25y5zEpRbQ/ZqwH522GocvLVXSZF+OW02mZoHiFwpE
axTS9cFKWJD9yMJg2kzMoBbuhah4qOu3lxPLZmVkL8Z9D6cHMexo1TSjuH1e2xBJ
ke2pU/OalXVhyoKZJlr7IBL5ZHg0VqhkujAwrQhYIBt1bhOqGYjycUyCjmSa3nID
vCTKAopqXyGpp0xrRZYC/sS2iy+YkZ6NnKrufJ/q/eGhtsaytXE62Hnt/aT/13gz
xba/NRbiP4z8LKCCveESV7wQhG50xVbXx2IP2P8VNagyyPHYqT/wXjezv0c7ZSKl
JmQ/9OjSMPMWNV5Nl1yvTPphqKHQsFRBcdcMTAVKcQpABI79+6u3sy8olTsrzhGB
AnVmC3CJZmORzlb/+yzuYOVE3GRONA7b9aL9YowLCsRLhcoLzgRzjWOps465Qx3s
Tq/gPH9Od8k0PQXPIfacKf9wk2jMkljfsZleTMipaoD/u7lzH+VKEDA/DkHuP4+F
IT0O5D1Po3SiZF/OyeDQBYSFjJbbaEGTI2VFKmntBK8XzzOBpcEq0xVfXMhAWPca
cprTxKE9VkmJAqVmZfG/JSB/ZqTYG92jOKPEfkJ4p0fDSJ1LxzNb3WzpzIBwX84P
c0JCOT2nehnBYqJkgcIiYZ9nTIE5pFfTptryvXYdePVVDmo5RsZuOf/rWZRbaYL9
Qum5wp9vSES5MWgVoPwY1MHG0x9FpJ9MybBOArOg43yW4CZJ5KvZ+yHjh4c3itK7
L7akC6XxoLmFFF9mT+NBJ/mlIQtqkBZZIAmG3uBsWZWi+TlqLTxBEIUAvaW4PIgO
2WAPpfVCiTiCA3he0GmSLJbHpAVZdj1QDdykIYjDqhw8fRSdsIcQnV5eQ42DxdS0
1R5OzksH6YxdGKNWrPPW07MFsBABKYVqRd21Zs7jNGWUWDDEJNAR4oSjA9ZITU7T
HJmicOzge0dKiOdvpOFncEsW5rTjQtRyhcG3TP/ykUpB0K/gPZTN6mX0JufjuLRK
pC+n3fIHuyIkY0bF9qCkosaSN0dUoHqqGpBUXcQ/ytDXIhHZ+9KmWr6p79GH0eSi
soTiV+3duQPcjX+IrqLqHdM1hwbH31uIQ605Zjub9VQk4105JGli/1ArtENXmvnO
YZizPgp6QHHnHO/JHdlYNnivD4nFpoIBhD1SBRZFBTxS0tSLBkGhdzi7qdc6x6M/
Yxi3WshyiZ9NCCvwLtxnJbFD4xRzQ8nSvj8xDLw18Sf0u1w/6z7vf7SCbOsXFRoK
ppZ8rYPrs1IBdvU5LhJnAq0KP7rvMq3fSJgjVG2cu0doSkwaTG8uVlE5TdHAuCW4
pcigrE0q09ij+PJinPuh7B3nvmzPFXCNmtCZbUApjAQ9HssNkdfygOgbDRcdWHj+
MIFfQHtglpz6VT56qz8sKau+yFUQRsF2lQ83D9y4vgYOBCbSfB/gNR+YD67nJ0w1
Iylx48McDj+7W2I8l7xMU/tgTudO9a5WhD6Bp6TlHko0iWDkmmBkavGiSR8C8JKB
nGYViuYD3cXhtthq3KN+t2a8XQhd4nEM4rKe1MHrM/b8NWet9uniQYOX84PP39ON
B1EFRxMcTgBgd2YIOsdnKBccuayGIZqV8PL/PQcxSJPXka/SjAhV9gQDQrPQu5RY
RBoN8ktVUhaRMX1WzcYyuvBPIsRVGrND0WbM1PXpiDXQWHr22L7XWI22rZpfGJSx
nGr5A+Xn1PRe0QNNZymKZ42jwymW7VjJYoC/cLAhgTXtiPS72xYX/3UTlCshATey
WKhvl7+TUUd5Uec3tKH0rcuhj9xJbraw3v9qeLLh+5oGl1tFRPGL298oBCdxnXRi
IjWclti0uawv1Jxo83K27QMy7ioZmYGVl2oPzzuIOrL36bJNhVE7TqhcmUNa4XuB
xoDlkZSxl2gaPLHgQWhlWhtLBZ6t2zrb4/AV8Lt89M7TZqXiX2KlaPwv0thS/b+m
1DJRTmTdnMimnS1KYzHaIVJFhOaoo7rc1/i+r9QFW5yctH/INGvil7Iw39jFH3Jo
zBHScVApdnD96sm3OjWQyDp16fKxoyZDGJZfoeucY0gAECWlX3ziQYIohq5l6Jte
Ro470vB0qQLQTyZqQMjubDAhuKW3TszvDXooIPnWhX29MUbRlF1wzUr52gMExBQp
mGMpDL0Yp/LLxQ9a5PLYwrTKUdndMRzykJzaD9QkD+QomWMTxu36K6v0NsNmIrmr
wbObEKHUaqR3/9e4ZQrxcDnJMtfFEM3hO4xp+wSFvhaRTfwtrueTe+R19G1SNqbO
xdVB7bLueXFWmvEl78ln4wB0WJB6MMg/1sifAHiyVYnvK2qqXcRSYjaCnlJTOwN2
rAvr7g5u5sCK2ZF8BPn55PS5K7RX7wPO4U+3c5EJflJ6vq3EX5vC8dnBSrzwnQaJ
4gpnkzge7EuhOkbf9L7Xvk57AiekYL6gr9D8hjoFfYGo3U3TQi8WtDKjWhcatX2r
ziTjoCOe3elCE5rOuRJEHvW/As3LXxTlcGUetyXxdNAaWBIS7b4H8NcGD6bZAqmV
3iJ2/neStLZ4WrkPXsgMI+ugm/ySdSPZ6YfXaxk9Ofi6A4H7fpoHiPapMZfbX2vx
xLPv+8BqxZerBAnOOYTaRDoA9O6JAKgXBOhUNR3k94tplo9LZk3OU2M8fBOw1nCy
IYOfl5XaFoOybG5UC0rNE/4TxQJs+gm/NbQD/2Wmub7Bo4WDbztdPy9dBfrnQciS
ZIOZt6/Os52IfA3aUR2MBWJIayK8JXxVHwIAtpeTM7qsUDp4fhDATNhvYK3ga/ih
Kwv3+jLRnSKmM/oL3nnAUMEz+G104vEqIBOFRJBIAYRiXNoVXnhKunKs5WLE4MIH
/Y5RAidW/dOmW87iIUVPXEzEBYNr0DQsxMgjGBmb4Ms0v89tIKLnFVeyaHf3fGq/
c077ctLevMCeUO/qdwAEDD5qw3QLcNjAVBAfJGSVt6xn9CK8aQwX9Ibq46NbJ9Al
9xqTuMloWJ4wYmtRhuSGZN2ZBcMramBX0fH/eZPYDMsnQrYkzF8t7wkM9EXG5g0p
E/NrePXKxzg1kAoQr51h1mdaUILSlCaRd2W5DNH1Z7T4Zx8qcLvatgaYxkA6VF6n
WZgmFJ00606OIO/U7uOu9hTVh4AgogrlPKFPvD/nRqP3ztVispwYyGTXhMIIFA+B
C0zdBQNaCglLpiXFBzWOA4jKP4dN/8VHSePSq9uFVnU8afgWtlucwucW6WTIlQcV
UsXhXy2/umBiyNtTprCxCDE/a/e6bXL2Xdkm6kdN/X2pzXcWvG0mInQm1seqz7ZE
42aDRVrFhRERyhvYYCl5nFIgMu4i+WYtYXptNQHfKW/DeCeBSPkd6wrdFH/mdQP/
T+P/nBcldRfon432zMCdnHVu85rEgWDBVic5CWUcy5xGrBkq+J+wdJHXUxNl+0pk
aXqGOZIMHFh6xVLK7qyPRmlhNX4mI5g3ce6m0HOvWnOkpbvKBLZ/prPuq1rg0XyV
+IaW53t961hhB+4n6Mjn81mT8DiEZENo4EgJpErNL7PK1pHguPp6bGXpcDeS3mx9
BadsQ2+yvOWXq4uAD/ETJJeRe2JLfWNljgPm+5yX2RjmWI+jNSie7rLbQOUBbtmv
tX/BsugUvUCA1gi7uRRoHXKqBy7WN5vhkgoxIsNtmM/0/0OH5LU7jkNqDOI5bUmT
dgpL8d8EbW5a/vAJeDSaLJvOtX1wZdXZ/DYLyaInI35B1riUOtIB9hAluzoh4aGd
MlcHiUv5K6YE5L4cqVSjQ1Gm88XbOuB7pYZDBRrGUNNhlP9L/dgyQqgfcYTKTuCR
5wjarZFIgZvF0CSYBA6X8dqBFf56hDVjy6bmM7TCwM6K/hmkS0qO0erF4qwNCcMN
neOQe6K4WU2OcCZpBGJ9Ec924Mj3X8V8RJupT/k/godRt0BwG4JdqJfcvJqQyTcC
jCRFTwHIHGqa8PvnwWDTodJ/JixRPHuaMGS0s/02f68BNXc7iz3XzxPKDk5EONkG
v9TO+5NwkiWlA9UQmEtVmoSO0/oTXP7jV5aVecgo8INZjlr2sEv2aPXB2a0xZpie
SjBeG8v3h8PeTqPerOWUlqH9QTJicl+WRbqP2YdTmjEoYmwP6PcuG0XYL+qxuyDG
wmmZSPcs7LyhM8vNMGQOqqjtdGB3jgyzO48tUh9+jEo3vU6XxOwjfyI7lkOXwHTD
+ECJXk1nqr7NOzE0aiwxmAwnZEUfgJ5yitXi8CGGJV1KZjskxCd5vcBreIbX9Ztk
YPjnv803GP0b6PR4+e0ldnkOoPT3DgXYhMFMIMOghJltERVgINtZcYEGUh41x628
OHMbJ0iqb2jZB5QgSrOzXc7JkN2OyqkA7YXvQdw9Ij+XXjn3TlnN74CKijgrsTIK
JmZIT1ZovUS/4I0vLQ41HMqApwJ7uyQ6lN16DjHAfGpmJxLX2mvijyTGJF6SI3Sd
tkaebTfnbK7O4a2h2EVt7q/ZAoYLIC5ttYyMXAJOO03gXVXberO7I/nR/wGxYXA2
olPzLWJeLoc4svv5UItAz/EPHXR74p07v5swi1rWGsYiYEpifpiYOC2xUYDzhix5
DDMRPajoS/UxLZW1HRgUA2Pd56VdjPs1ScjPcEmBd7KSWwFNJrGgx5VKgVoVKiH0
X7OSjioavCrgxB0q+sSGZ1WnSeMq8nz5vj+IuA/QQn7TI5P9DuiFYHRJ2jOvw9T3
Auqk3kn5JPYOV01O3oxfO1LEKLijx8hKg9+RTZa4jXUGC/mHjfZA0wNeXWf+Jyph
Gr1FYb+AGHFGgghrDzZ2+rWRLwajL88ZxgMxg4tKHOKA9hIhVKywzBuKzaIUQBGT
u72dzy9EXmN48hjrnuDOokzIXSYh1Re4P/l12dGnQcIeohKVd+BD7mW7TerTPcQL
cMT2CpF9YbcFYOkzOGlc6NTI+zoOxM6pxNKr3PftToJAo/4J1NAu5z+pvutxLdB2
LxB1nVy2ajJ9+DhRTMbwHm50sIuy+i+c7cybW4xwUQgvQb5BIy8IC/FOpa3v5R3n
rjdrgYVrgAW/6M53lCm8AWVKxYkmNpfbtDdA/TwVijToyySAzTmLg1sUxnI40UcE
Q6PzZTu/dplA2gwtBVINoxtDxfieLNul5YyzBU4z60uxHtTLOG462SB2GVAAvAtE
gQ+OTbHFZr/OPA9J8o3VwqVIYwayN5uAIP0omor0oGOS0VsXn/nrYHLuR8e4oKYj
ZoX8eNNBjwPy1S5bPaHMW43soANWPyFzuU0sK1KOqBReEKkRmnfAFzvBgCiksyKy
ohoElY10n1iR8SaFbGJX7QrLY1C/jCNvGyd4lJQBI294ZNGs8vO6uI3HnSKxmrJJ
OeP/yEOw0ctdXeSA5sLiKK9KQNRzgzbFvV711XO/NdJyk3Rt2MaWnuVn2r2VqoOV
tvyUVZWMjPxjKmzw3T64ClkqmBF+aLaWCKLLL3oXi6S9NzqxZqXj4ezQWlKHsXTs
Obo1lXzBtYeBBnzBMVo8VBgNqlEgggQXaqQ+wnMlIQberAjFNg3U1cNHyZ4Bw9WK
VAz2aLYaoHZxN2pD8qBBJLFFIRXVMf9D73/DCuFhdjJ93x2SUZ2ILx8PQnC4suzJ
/kzmgwZhIlbix04aVw+TDGrfdtcZgN29dzaWrLqnXNKYAgjVZgxqUhDr/mhPBrwX
UbKxDQxaxZKcrTdBHhT1mcr37JhuGR9mzKfFSbBG/3l5vw0JLo/zBzNQsvtEZa9W
4S+tI4Bu750dZ6y//YITxCXrkVeGrlfj/CSzPnE1+yO8Au/TrtOdul1YYFoi91Ls
9J12oNDKwwt8IHfXV7SOtQTvy8qPbLNJpTTxmdO9kr5KWWlm54N/FdkfKawaV6Be
AjfM/YH+a+hSpMFxfo2NO2pDeIfA2IHCacom+XKS4UAcFTud7LJi4I/PFNdmD2yX
DAIX/mJQFoZxfky6b6AXZWlqsmAB9qaXceL2tGgkzmx6/ylxE2Cg0WUPowxThbhx
ofpe2ltqqZXViqAuKrTVn2+DuZpmCwpEjT9nZn0E9Vj+xsN4LvnwbS1g8hfm2fyw
YiXDwOxO1HCftfrprfV5BEYkorrSglMkjQlZWws4oSxVM1uf1tTNAQVtGifKKnQK
9XROH3eeLjd2A9EJiTjSrQ5WNv3kPlsTGfPp6uyN0oGWvpnyaxddIUBW9F+iD4ty
aUQHpcZfucvhsCIF6gYxv3gafcxE8gjhB/c7qQ4ACsP8Dy4kONvyWsUVB9u3m6xQ
oKHpmLaodZahKbAzwx44ARK6fAF+6bE8B0Vtutx5p1EdQLEWpzaH/cquOum6igx/
F3X8ug/Q2gvHmLQtUbCTTGYIYsOBqlB/NSG2CyGaPMHo+4/oZGhtQE2HEMJH3dfY
sxvB9fbiKq4QvYgqKtO6mDxLJPv1R+gvXiON+1mGY02+/S3ar/y2swv24p6hDq3u
OH2v9plxxrKNsNaImv5yXFseYXm5jzPjzv4kDr6tYAABsUwYpM7sOEN7693Zu9a2
ZaKdyTDo5Xe3MygkoKZQBzfkhxDH6urs4pzq0KAstUqjBYYvbTnHFRk8zblhkryw
F6Xav9RJubM9lxmbFF7Ql8pnzdMDVjQuv0CU9lJXaHJHIzO2M8effxL5u8FDdmnT
9Lhegl/owMnCI1CUT9/a+MLuNuYa+OGPiOwn5jFlaY2TsYjVtlvsPM19qDqknz+g
vHQdxWfWkqogSOcKhCTuomfeRKMJyWuTzl6/re65nA/3NHpRXREVnJJ5n6WA+3FD
2mNCESB19sskurcncZOoh6Ef1GKWzVsAQM+KXuRZnPNa/FEV25ExXSKAHHDOJI0F
G9TxXWc9DAP8z4tuLTbfvx7XK9KpBJwttHiZDWP+EwMp7gXsp3b4tgg4N67lkOl9
K4INIGSiEwy6TZ66Y/lI1jJB0Z4sNDCSTHMCy2PqsDh6tuu2b0NTMQBxcFmG1kXH
7ULGW1gsX+TQXWI4C/USofIb3j64I/vI4FAb8aRYHPUCG6FI0GKNEjrPrqKj/FHw
y6+V9YIoAF1TlaUAExeqqKN0ZhGGcCCg/7blGNiHKjuu2CMj6gK9FFz6hp8XXTid
jEovoTV2OG2ZiaswFLWY5jzLQXymDkxLJr6b9vx1YHK8/90/W7gL0os8fZHUzGmQ
HHFEyA9+Y6gcKxXMnY+qPrbDzdVni2OlKB+RSfTCFpaio5dskRqTlPyyDL8Mf/tT
NxXHRwuu1IO09zgsDSPO39aG5gp6sZrYq5W4Wu8G9yxfkPTmioD8M8JEskS6/Nvp
yaaWIdmdAmBbvP+Gj2tQF694h1SqKuBzYREfb3dOfWBX69v1Tpbhmx/oo1mujmlw
YX+L71qe1Scw48MdTFqTUiETlYvG89BV3O21ovZu4aQehEACiVG64Nz+0JuDcUve
ssLGmeCMLcpgi2FWXBbHjA+nZW/7kiAUiGsRsX9LRvvhiHxHYIuR+Qy57pPV8Rvu
1FR/gRpsAqlh15lzHUAK0rmZVegDCFIOg4MJArIhL+OwAHdsG9OxzFTpPxdxGKmz
ohRlQszuQpZ1qdVlWEsT8NfVTJAJMc2Bmzc2qVN0Gmx2VZ5iGRpM70pyVKF66NvF
mPLBp09HQo9+tqm4VOz3EI3IapzTJCG/T5vmHwqaOOpcrntGVdf5O9qpHtHUgde/
Be3uvPNLoyKaP0JcTKHgycPT3ao1zEUnVxNBR6oKi1iJA0UlgWZVjlEKEOOVOCA0
69l4DbUq9I7u007sdBSeqDRpBs4p/Udzzh1N7ZcuDbKw4vdySCK5BVE+kB0Fw7HQ
8u9VdjLpEgoXy41OGiDMrQkz8k/NoxE3FdCwvXC9IeXsKYziLl9cxOsFbSs1rOVA
GRJYoEMRxWWK8rL3HrPF+ttcJ/CxcjgLiMxVeZK6YGqVi0pqVyjv4wRgJEz8c3Lq
7lrGaHjJNWyHox27eDtEocNIwuoRmAPG0+JeTN+h4oChuc5Eu+ACM3MAE7rrSxzQ
EACl4L0D17tF7jAO2T/AvDTyCRKQEpnzKXaxoWVBUqwv+CrgAliRiCfPw0IMANc2
g5diY7dg3sLRUhb2/kKK6OjvJ3w8C7zDQ23g4XnAG7HVY0ahkdyn17YbxXS7aT3s
RfHKc22oG/UszEl88hWS+ijgEGhH16K71v9rjzztU9VW0GSo5QoRK2T1IskQQ0Hk
9mkq3ERuoUsbLSe2mlV+ykb9NusyXqhEe0ugyNJlNf9Oulrj4ZKr+rmjdOvktDOk
i5FHBginXMHJk+Iv5PXx8qT3cYERgFPTXXFLT9RHo5aaLL11TBcKwf+Ea5hf5kqi
H2PPVST/mKTbxHuHwRJmKnLFq4RlCeAP/OXzL+RPWxSBgaYVWgqh0Nyd4Ik0FGCL
710m1FyOiCl4C5/0OEY5RzbId6+Fd0DYEyx2sf67z0hHmdIbZNgjAXMHD78k61I1
KNfsS4pLNvMIayf3aaHfy0Dvw/rB9d/JiWlP9cq1M4acaQGO5vnGVJIfug5LOkWI
9RaMKgEIoYM7EmjqKd9ajSS+M7zcNZQzNhqjm5w4pZbHxt8YVWALSyFHR9XzFZUS
dMrBwC6YJpNIw8++TyHGKl2KxISUIoZWnrOodkJu31Adkwuwaogfm9ILMYvApZX8
qSnZSmUq7wAajAbfIc8W+LXYGa9iiZOqyQOOqQUogm/hvuhzNjJmCqF+CR0uXrQY
R0mfrKc6MIE/HAPJeuoFFSL+WPmW3rIeg9lJXriOKk37AAl4wLJHvtOsP6osHtHs
wF0WuIda2iVj+kG7SG2VXfKQm0/Py6vEw8HdvTsDdPD7Ww3Y2PmU4ChzOjwrfwVv
cC6eUF+os9GvW4HlFr+K1HGmHccaeEj1SL/4nsFISYplgDPoTycRXATNQEpD9mIi
3EJGBZvRBMD6m0DlUoCzPOQfKfe7IdMTyd+WwBMPN+VG37JxN6IUrm8FdjtXej0r
M7qDyRQwxlzG3AjjNTFBV+kI9roEvLUzIkN6Xel8DP4nVwql1trtUi1271l6yypH
vIdGv8octSgAL7Vsn1NrGLobz6rwtN159jmgZZYuMTouxqtBz7Szl0OqkO6/Hb8/
WvEjqJLeHAocc9SW7Y3tIe6j7gm/30jHvVbUVM7wb3t87eeCdM7nkVm9mEGFGOgu
l5HkhX0OOsylOzyHpNslWPCHMSR4cwJNZSskfS6oweiyqz3L4jfNyFGKZSq4rF8c
XiCTS2mAUfzVYoZtlF7FBMB5LvShSN2IvaTYzOTDpUp3WxUVVBFUrlVZrub5/1Xg
TbLh3Be1dYzFN/JRi0MFQvwmiW/5ABVLTrelCW1EwyGHlVL2l992yirDmdxpnN5B
USviZEAlepNwDYyFRS3iKCTv8X1a1JiAfR3Yiul/ZO66KDE0dsWmHkpvMchwvAP3
Mp6x/WV/Ozr5zWg11O9Zrmi0FAFTyZ7BZgrSOui9W4JBHxAH1gaQ2YO30YR6mR4j
f3R42ISsYs91IK/tWT/zc4F+REs2ckQ1gbLnmaXqkdXjzpmUC1IKCDSOfV2toCqR
dgMS3rUTN/VAMoQ9NwHnPTIXjE3Dd3oVOAPqKf3IUUESJpdEcx0UjmZvmeG1T9vJ
TBULeVgPYXLOJD5ubFlC0JO4vEvueYdKJaZ2sszviFYU56tJgwO9X1NkfYDNaKIN
o9Lno4Fppu2Itw4oNLtnXjnsvbpArb+AR2pC9s/xRKg/7mLIhYhQPMe0QLWUKTJ4
f/ggU5T/G8yBCD2PH2x3o/ugjpL0CrQp0XA7dHZbcEBUbNNCVzfQbj5w3dPh/iep
g39+8ySg51KrJbEaimDT5Pi6APFGBjbDqMUZVFwBW2z01CPryZ9ea2obzaQ+vK5c
11aCEDbyoiT0yJ6Dm08dp6+YoU+874Ipf5br1PuTIqVewbmHK1XPsWKqNv7OCjM2
+1szyK9xA/miLGRL+M93exZFs672G+mrmNa6G9POHJvQlaZpUieTY1TB8psyY26F
SmHBDvuo0u2pFMFT6H8fbUl2InozPvDDw4/iRcLmtBeTUZqWrhZEOWSErsD6WUjH
fgt1QllBUi3HmURoOYmomc4/QWIvNOZy9J1Pjm5sAWsbDaSCkd3jaIILyaJBrAEp
MoK8NG3+ATY2YuYqG47w6ZtWMlnXf+I1G05A5UedVjEtJX3H2HlRI6MzU3TYNZy6
e9c50ylq4jGL+Q5lEnUHNmjUtaq9RI79SqJ8I9NxR6sKoCoe7wAe6cWLoYq6P88s
Yn5tYa301Gk4kNrpFxPyoFK+ceVSynY++qYTTz9A6abwsRlZTr79OSzaclu2lsPn
ClKER510aQphO/tj411HEncZnNYqNqiaFMmxiEsXC0XpjwhTI0U5/2XYKQF4xT6z
029msKlUapuWwPvF9XYjEbJd9vVx0mAb/boGjGtCGutcmjHxo5fKAUmHCl7xrsVN
1ZW0iWBrcegTTs2gXRBD5YVAadHqWsBziglLMz5vMXewOR8XCpGZhsQfSnskEAk6
KhQr6wvwq1KXaEnFFmCicRCXZlptbh2UAb7P3Vans0XUX9Zbf4oHQtVwynabejXb
aVo2u48jG3dyUve4XQqxUHhGV7mk//nE4pRtRBjtA4s0vMnBg66lxJUFgK4GNjgJ
Dt9a/ZeasiqLKcpGHfFlvr7/MVLRevB8dVDsjD6vs4Niy1ZpcvS2N9jLsLsTxRM1
fLog0wViDj7bbe1WnltxtgJGWTMX/yM0/yObShszlhmQZ+GEV+LRDhJXB6vZtfVk
48np2eLIrcguA3klaQWqADpI9I/5VGndVPfOlIuKr1tFqn+92QbSeD+YyR6oD+1S
APeYa1m76hrdpDnwNaXpAkT3QSBTDJp5A4S+DT/xoip1LDPoYZ4xpdDzksIfOjlX
wek23w/tpiRMPYeVUyHbBT52FLTqs60LbqJPIIJimMtbnMq857DmTB2z9SX604L+
wfiQV7zFNExXFCBt6hTK2fjlZMM3lH2/J5QHwiu+8LKQoutRKQYZXZS9tdSpb/eQ
FcWB0YomDWccrINe9pcL6QYsZswaiYTC749VGHN3L6skBFZlgBiY8Hbf6Oiyjv/m
R5uLDrD6YUCnqUNk92ajeJ9UaoHTPxJ5M8seUe+zxA/F+AibFFsLxpFAzzvIKY4I
caVyDnrrkaPGOh809nsvrCadE+0VKWgmutkNJnGYUfr8i9fcT0vYiBKagWngtVpD
d9is7KVUcGq0PB3ADRbaNErEbTBBCJQua4liaEo977oDChY1CwMq96qhqYDuDX6H
NqKp2C40ZUy9qHkyOep+tkkCMVBi/MfnrsFrWyg1y0zjr8voQ4Wz5pokE5a9paE/
uGWBvT/rYzhvp1+lU3frEWN148ccMudFRAA4fQu3/J2RM6K68wqIDRS75c3ZOCpy
AWVmahHW3x0OLenM9hm3NXS+H59p4cPP18EHlyZRx4CyM5o0/y9rDwbNGxMpDNUq
NRmmbIrFG0e9NU3ztmwA9WD/vGHyjjP8FH80Bo9YzNZt6w28J2o9sMGdlU5CCzbz
EiLveFUxgF5zuGfTeugLlkt2XHBb2GJdaN6vSEjni1a+ifGnrEcvBYFN7IlCYf8A
ppNe0VheQlYMBbtF0p7XdmZYXsZdOpGw0GT6Bs9s/mR0FZObmWVhTa+BI5nlXbNs
v1+o7NCE6SFzZhfIXo5W04NhusfWSJ3PSJw8FKQIrICO8MB81UGF5SnmflTuVaxM
Ypq5jnUVxE+WFiVFDSUPkwLz4idKVGF2+fWfQpn1Zwd1l+foAk4yQ2oKEcsen7An
i2AYtocT3slNH5b7eCeQKOS9FF2d701JRE9E9iF06DN/9U3G/H40YMNhAMAOjKaj
CHGtnXqLr2HfohV2JE3YICCWwu561j/Af7Qbb9aqV/eOw6kojDv6mz1TMb/xzsx/
loMYbMM1SdqGoYdMc3aA3JiowNAlXfbkfH2DUwSoGX6fYnWIzzBG8A01BaZie/eH
bQPNFncj0KX6wgHJ+dm0MCDiKW19PAnEzsaHY1jGru8emlXPLDHRUVt8DTEaEaOi
4PK6g/dy+rlr57cuqH4WcsvClRyEUDMO89Za7VVqmee0ghfrcTvqsAMTD04fq5BF
NWRja448W8i8Yo84M2Wee6UMrYEk9f/2EWS1xE3kZxi8br8gaEhtRZf/2tpr/w5X
Vj4AdBNwAKjM5wST218o/AE6gpSoo3ECiIrBYpWdIPXXTbbxuJGCW1/CYuPsiJ75
D498ImcJw0t0kzknRHnOI1hKrwwYsE8FiRWuPV5FSZMHxZZ/CXNHiYsqZPp/Ifj7
kIk81Tnowb4mOGd0uOeBGlXyZgMePX9WwAtyzoySfdFknDMhqxo6+M7ON8HIP8R7
I5Wkam0aHelMKiM1RL8CUTnQgoSoIqYPVo6TNZmDBH8hmgUwaRAhR9n/5oy4deVa
2+N6X8zG+D1ejWqscKaWoqKDP6TtFZKBnR31fZrsL4Wh6Hyg6jVOUSmSTnYbkGce
9bIjeZr0kOfbtVQB9+nbxLxIo6vzreVfQrfalvg/lAboPU1QJHouXs/evzpG0+0e
VKoxUfVgzbZX5WgKc8KB1N8MMWaWuvR4QPIVBCenQQJJInftLNtMvBC1A77/BvyZ
EW2xNYMWbgb/hDbvFDTCusvQnLi7UiuIBfUKMHd9CLg5NoCxQ0CyetHM95OBlCY7
Pk4rt99v3qMnLKSmMv/pHgeIp41+WqBg3Gw0CkmMTFQQpPvIBNLk01u0MEOlVmCT
C75M0bkDkTBYCIEzPb5W1o/xFOJFiiwBCs1T6PjYerGO3Ij8CHTjCRghFMvbJewJ
paTtl4iRKYpnSRU83yu6SFDwzmFKkKKKDzz+BgiVJHHldX0DBVqVRreP+5cxl4Q+
w/BXTJ92dfwZ13eOebqNavMFv7KajSoK/jbwqgqqhGgUNtBCwZNdtf7uQ9ruwCg8
d4Fh+A/Msyqn80K/WJY+cSc/lsUA8xmgstFMTtswL8Uz1TbC1o5Vvk6c5XH28UAw
c9z1Pd31GM0TTaFnUNyvhONbDGmlM1593oyLb8wDcgReX+UpKeLb7wzBlbRHK515
NO/HkIKut7eJAzA3XwuhSyZTLtRG9tZyyJastZASQ8mCoPoVJMWLK2VNUvB9391f
yhabbCVFodIKvsWCGUGG5xvNKlPQ5l1u8stTHlYVcijAgytcf1fpyd+l3VrtuHLd
ch1ZRYfAinDoEVvot9B21dc0nSGFLcIzhytnzCyHMhzYMaz3WdDIerAhxZQf0edQ
lKtDKb5yeZ1RP4hWxzFc3b45zmbZsr38eMK7XV2zQ2ubajpCovEmqZgHS71O2jm5
doFyaUfT9ywqatnsZmGS0Br6fWv4e+6fP13rQiGYz8Qv6fxWa3jlhOpVhkX5lpmr
VMJpB1/xDAuwRrtB6x+cO+wCx1Gb5VWZhekBU0zX73i01FSoQPNftdEdmUR1VkZo
/SrUU7uAIVjw+fgplw4zPvGPWGRBILBpXo6wIj//iV/DcrFTr4vs2PGzMlmXiZSY
FTs1g31jTF0Zco1OHq1d/2CmfzWIjL1DQDvNaoIizgLiGGpMf27A/+PgOqufpCGv
Bl+EFXzUUzmzECFQQ3CvdPCvIUtEll5qSxV8qTrx/K0TVYfJCZ6+DGpqI96AR9uM
keArZEtYz4rTM3ZQZt3zY2ATQTY9nWMgAFV6p3XjCJXXsAW66XvpJq0JsqJ1bJNT
fUFD0g4Y1d8Zxf4nnerm4sXqaMZGV8uKdImNXE1VNDkpZrg4UQvmug0eqhB46LYp
F+sv6jetcxZW6SO+jiZow7RX+zxmLihnOILV24CKiCw/ZfO179wOkSUoHZhwQnHx
Fu9KOOiW2GQnL5nylJeyAHHuxxoP5RGhzVSWMNnEcOU7+j1eJ57uSzv48peumeZ5
00t8DqPrz1efaPQKfenh6XbqsWiPB8TWd1g2E/Gm9qemQlEWuKsW/R12268fTLIM
WM7UXQvyQ31WNnxr8O24dwt1ZYPgyl5gnnLVhF/wz1deKMrorl1q/fOTjnL//fv/
rLybD5euqPM7sHgPr0NNloLGJlEIEUK6Jbh6L5uhDwCIUkIa7XZML/YZ5kxOZ8mb
DeP7KlNde6+XiUV9d0vhw7PDHKu4CDN5Oj/rWS49levJTztLi6lZWk9eWlEOxfEQ
f4DzPZhDOKAQ7sio90uKrMGsqeGC/b/akp6JbBeDqs6hEEnPoM9k2pARhNwluUX6
vQiCvkCk1ABTpK/o5b1Q4tlCrGnGemLOy3+NfJiIz1fzOsZk9ln+KjMoyg0Cxmx9
oRkhlDorhB6z4+7Na0DqE1vGE0dJuDpwRur66kGyQ369roK2iQ4ZV8bHdCIMKtJ3
n720tU5XOHGDjxkQnoC7e32UvlyPR2Nnu5TtM5YtjRl/YfuMQG63iAbAfNLinqmT
XSfSUTJijGiXMuk1Bew2roNZWk3KSrZ/+OdbC62/HcEo4fJ6VrJF18xX0W1OQEz6
7RXCwr6gZhloeINtpLYaw/Q/u8dXlZJ0D9m1LrZRqiX/0Prq/imebLN7WkANOR2I
P5F0ur60/98rD1HzAav6aChsT0stM4iG4pto176OsOGak1iocgt5WLA3aOJPZd3d
PzbQsg8gych2QySyOqL4U8Ux1rgrDGF6xWNFqUnNnPE1WuDOkg8MWCLm5ZRhxyge
TXn166Ws4vnrKA0WMSWhd6DW7InaqNJyonMCT61XCwEJaKpgbjIvoXLpoCH9vBkF
SD7lzoZoWsMN717FAExn6mfSOeU24yJ1CJdepH7IKFDPVArDOG4WemqEW96BFe9A
zs8yYjeS7PvtvfrLoGc2R3gkRzS295JM60gylOwCuC1PLNfRQvYMnm0WNOr5qyIq
san1jF+/AUN6wJhXk84UOaXgF5yMkoT/a29MD+GMzGki1a8DiVUPERNK7q0Bjhvr
cweCKCWYclFiYJQOF/3mqmXBivtX1HA1wq8MzhCyUq0w12RmFtNYH2hQ1i+X2nXG
aNlqDl3TDvEIcCybfMQvmnhAEPPPZQl37oXMd+yzGLeXZIX7OeIWsdOREgftzgQy
jb/uqBKE1AkX4tK2ueUPK8ucHG6hN9gs57FmVrnoQqHUNJI03H6mfJwndK8qbzYn
tW1E1M97BIcznWlQJMGNObJCDul0/osYt+JiC72baeiymtAhOLwgeVbekxxTMtVv
rHkavqh+W0cFDNyG6Q3TF8kXl9iaDTbQTTt3zQcZdUL/HvqxTfxBSU+w0Ob0Qx+u
yfIOIQpcxeHq+1RJuE9ixBa9arKkdPcdNODdPQNRrIyppfYgRXFEVe1M37X5irXd
EXKmBPXUTxTESXxiJszLxATUvidJliLfdEDXxYAtvudoLw2dZnnm1wXNA6aYjqIm
VeRrxRBEoXQd/CCwqc9K18dZ6Czt6CT0ok1vNQS5iHuMBSzb93SQ90q67rZnwqHZ
ALgo7WkZnYSqhqZ2Ecps87UzJgwZ1l7nr74TUw28YeF0gjTie+wwC4f4piAAdH/P
FCvnP6YU8UiZIrdgczIJFDhhINsIU67n6Tfbhauah6vxx9t3mJBtRqrCB3s+onms
6tNJB3ICl2d0ZQRuwVpQEPzjOSAUzMpaLV3dSk48DKWXkS4vlAQic2FnUUEmhiC9
reDMvkt6l6KV2CpwY6eSMUprj45TPwdPFybxZqFYmdy0rvIY/N1+uDKuv6VglNsB
ZkT5d0zARcOoZD33gj4aEZfNxFpowgHLSpcmSNhTpyZFfj6/GImdeF+QOScimJ5M
LljjVV09JfeGnxI7gj1+AiYPFCbOH8Vs1GCkF412o8EFGHQH+I+LYpUhy04Qpe7o
wLJMwUVHvNLNJzQ/4rRx3IFa+gNobgacXfvMDUevWVkA6BaAqGFkCe9hWdPMxwzB
6HkT/ycl0Yol8l40wW6OcLHfdVB5NyrEk1pfJeQbkEHAiu5p8Q2aWLfmCCR9J+f0
/Ys2oh82ZVLiClJWk36xeGuZbbpHJK4U1/Vf4Wd8L6AhftVjSi9o3/Q5TjppI/0v
lvGvr4iHitPlMY5fW+dPq+WSNh3/SXDsC1+PG8GzEcWv2NLfQ1kJgFMFx+KBxxs9
8Dcb2W3Wnsrlysx4Ee391dNBMX0gh4OCy+O7Nd08n3270JC6koZHJCZ+Xis1Wv6W
j665kcFJ9yeOEz4a1re5KFlw5GM0qjtMgkiueTHyM+RSjGiicCWiCyx9gtKbTrm8
wKorwoOnMrZXwBTzWvrPOO/KqDVUJmPQRDKUMlw/2t8uTrRX66dvQ4A2UpBAajvY
dwH3RlhQS7QWMOf2z29inqMUPMxY9vE3JjI1cK/T0KYYUadnC5uvHoFL31mtkwLT
fQGt9+RjuTEsTP0xm93TM+kYFYGE0cMIpk+7Gdr5UVCxls3NQJLQndB0AEZu0UJb
xRkjUcYO2PW4YJblJoZNOW69ry8BydshUdjBAJKl343MWCySGbRf0ftURqvtif1E
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
URPcrbiiGg+L8+lrIDjFLBmhFOonWmgQ1/S9mYSGBrzqfvdltwPRvTro5EKi9MBG
dun7v2LHeZGnP8lRMmYYn5/F7RKkYpygVvU35AV5EI4NPgB4yK9WvYMlnZAmd+Tg
zI2seP2D9gMkTaHPwbX9uhiQ1DQl/nhZ3dySGMIBMcVPSSzGOKwyFLkb6HsNeaIZ
SUCL554lMwmrAFikw/UIN6xMN/DzFukoRNgMsFxcJwFpt4KkYqo6otvR9CrWvb1M
BrhmMluG2ZpPIu5KgNL47btEq9P6ijWHn1A5PmkE21zMlmfP09O/T+XVHc/6++rd
hW31+6TtXG6WEn5ZEhynnA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9568 )
`pragma protect data_block
syYuND3qBi/+oDQ6Jywt5obskx1EQ3xifR595Rlw7QxiWZA+tPqVyoqp9S/yZxWX
0a0uAT0lvr5X/z6g589kLxkMrzieYhxtwX9gvYpD7sWXO7ZQgC+gQMUrUX7OBz0l
wE8nIBsdv0rCRYUnBObomfl+cX4nw05lNpeDiYyz+WwY1R9wQATJh6CuLu7hjpLa
RSxpfvUQMrRMvDgR875vgaYGk7Yp7Z8ySQx2swwYj9aiodPuaQsu/k2H3DUywP6m
3c7Pnyq3CW7H3pq7WwScwMcI7RMel1U58fVsMcD9SVjSDZLtf4QX826GTdeUvnmq
O86wfUai/kQpfii4eDQjsjudRthHrdWWEssYML1T47ZKPeQnNouNJAABM/kpb6tO
MOLrVU/2AM47mo8RAghixKsti7aPRerOdqjHTZV6WjaKTBVI0cPs8w1eSnXi+biN
jFW5+er9Oja80dW41F3ubox4XYYjK2Wjr7TEKvriXJVNeuWej37Sq4uR++CxuzQN
btPEYWvUUxcSbGcumlLFpoSeqktV5lJetZuksiS8VjnQvTJzcts79UM1LCXqU2cD
EVbpAngDAgzaAaisOC8PJgmNfKf9NIEYx/sIgX8D8ChIFylPToASmtEOCS0B344o
AuO5c3rJPTx0XoAlX8hlEyqxWvOXwUHi9qqHKRVGMxA9a1CgHejML8iX4Nlk5RlI
8EvBf/G3305IjUSgzAI9TxhD+SmXcM8+mKezO39LTEPIsrrtudCM5cOMRih5QY/a
zV6q1Rj4t848KhBuWZ9dZbiMeNSGMVeTgScPWRFDfJe7X01xNA1YUzmQV6e78/nO
9U53V74LYnRxtgQ8RNoXS/nHmOURtTGA3NzOEzYMtxgv8DaYWx2zRR2ZnbYwSxRe
iuuPWVUp9v3lp48+56krgYahtzBWva/v7RgVZQz7vjZPiOEiNRzvyu9wRdMXT1/X
Cxq4uJyLKET5nASG4AG/iz2ETbZuXjxgWgQ/SmpV0Egr324fPlcFqBLADoXgct4B
tFE1AsDaHojkbHZduTD2mAHyO6iuWAYmfGIAlwb+PaO3BmgKnrGft55qisj0ga+1
WfmLpSO/kAG7QZeUfXCE8msP986piJjyi+VpDvYvGKJGPrK+p+RCbCuYn4bn/Ulo
NI53/6XMmHxWFqNy4X9hJMPUKdnjz4UIKa0V7OdVdDnbWJ24osGjtiwVo8fFGKwl
yX85pt2hbxOMybcLL3lo+5rt5DmzbYtjVm6LI8P/lLVvAV/c+dZ/EZlmaphBF6nW
hqIOI0zY9g5rICbz3K1nM8cQpUIcn5kUvGKKtVF3s5YhBCfU0LHjTlsYAYN0BILp
SmwJ2sNohnxTySHSLsJePcAAxIByFRzoib870xxFklbWF8kGDnCR2Y3E51z6HrjJ
sioB594O2elnLx8QUn6sC66Vm/Z86vcTWPk/XqlJA0cafVFQckc9f+dzlLSuzoC6
ffNUXz/aVG4wekgnO78Rmi1BduwNo9sKDDWYxZXSGSbHmZtpXigdSJmofjQpwag3
sfarzLEjvNUSViTUYUqlGyGDGPAwXA/tz2szwM3tUv3HX8hIFDnQaQhlq6rbtq5G
rxw62X7vxjaoXDJcpLAwg2xgwlHZIuqQu/JXSSD2uKJg6gMVKkbz9qTWS/LYf/WP
IVAMgwTQhlk6OLPETQDMetx6TFhIi6LAK1HMZF2vS7EAt4OaBdCpMD8k034TRGO5
mlmj7zaixOwSwpLK1RMauLVPTJQ9f0BI12f2SxtRNSRBiGphuHQFayyzU4jHDT1e
7dU/glfdWNhuANhMJLSlJMAFZVdwxDvKGpbH4rO0Iv1UBgXiIBW4LgZCcC7cqpqu
PBqf9e0QmW0/IZBRjN1JwUeqCqlZMgtLFToTVJAC7YV8tXnQSMcfJZ/2rDXM+OaU
NV67zCM+P5wYWzzk7IjVbzxUypARepw2frdnQA6qwH7gFqXqnv793N2JcJFk/Etk
B8Y2jAHq/Cjuj4YbsGcxAV9yID6cCLFrWxewAi031JKjOi5PGU69uEkvvvcuszc9
LRdoKeljBFWicHSokSIVh3r2TMskrbroGVVAM4Li5khog8i6/8Tcbkf8d+i0JGQf
9TVeSCa1gczKJgSeFzZhlCnBVkF8MmUX7H/5XbX51fZn32tqhe4SzAwP/EIKjt37
ME+M0Z02bHYnMxS0ndvBw/7/OG65ZPy7dRc8U+CBQTfPJOss2wiAUmLb0MP2NUNj
U9/kjNuyibI0U19rVbCbVnVlSDcar73RCiedaSNlA/LNRg7M8WDbL1tYpdon5/ab
gSBuVUcJzTj8ch3gR04xwob2nmSLl4J7UdWswv29hugw4vR/7+BQZMRXHwmqf4Hu
oLkEnFRh9ekLEF0v7GedqdHp3O+4jI0O6nHOt2eykhXJ3a5thXJa+s0hT7YYg/s7
FgbMN8vuWfrGDZBy4B3rE06hTLnYNvkveGXKgeJE2PDU+aB/Pw3XKyLvxpePYnGa
bzQ/vg1kmA+w4HvZTa7ozHJsL9y7j6QcVVxdhmMdd9DAVTK7HGkkwezgrBt85HNm
XVCspa67HWsR6aUJp1VogLgbTyFsXcabYZqf9bl+ETyoWXGuPrj6dVPA2yN66dbw
9e+ys3/HBN+A72Sk5DWJ1+Kdrma/lgLvRMWqpi23SNlFDMjSWvA37SxIgZ2ouGVW
TNiM+K5Cl56kt9X2h5ujWI0Qb1uIjxTwSnTQFpIqjglvZbz3P5vemxBK9CX/U/p8
Dk+wOc7//Gho5X+2BibLUxkQHQ0E86ZAh5GJzAPwSalrr20g6GxQx5WdQwYZx9jG
Uw5H2myU0DGXjsjqLpowHXFB6rOfgQVKbGeGB2e6pDUoLFlqE0I6jJpIzwudO1p+
y1OAFLj0q3yJkyvJSRlPFDjQn2mKBF6czTZ9oP0PLLNEhGKCtgjmt6NWd8SHCLhd
M0irxd9cXM+RnKPCPqIsOvWaeMfHy0DwIJgdgxnxXLKp0L91RPfu4EtXpvs4oD3V
btjbpu2gI0PSbnnJl2Pz5HDrJHBrk6UpciCO9e+hZbCNlvZYmCp9mpIn0+uxIY21
tRJFDOZytnmCHFaSqy8S9xOE3jejfIzYr86jB6kclhvQmokpnvjOy3cR+N8ZpVBf
MSiKMUkWOe3wrl6tsP2QCxzzJXvhobVmk4PtyS4MMC2uLvOghnnXAyUCcJfxt26D
gOeqEoGKW6JUz+Bho5f05hbKA3Ym6LXMYXMi9vdHS2gSCvdazo33CeDZyeq0vqKK
Cl8e7vDaLz0kBiGlKko3WOvjg7OplpYR7bH3bcPZCF/PevK5x5AJqJMRxfRBJCrv
1kx7PgS8owmTU6Ruhv9p0CDBtxSK9phG7Lm1zrXzwBCYjD4O3lZCKwH/Fk838/XW
/enMIffmnMlGxzmciu7bF/PTAsJeeOM+hIZQFPL+oiqgmiNM4rEFBqkgz3Rgo8l9
vg1QBqm1VnluxAnpPGGgjFrhH2eHey+UoyYLthRA5P9XGyrUK6p2/VIEpVwLlNom
bwhvReUoiGCM+2BjYUkkZIViSlg5gl/a5MQsB4nTI5b72q3o1spUoQzygdR/nmuH
G5kBlEfdl/yHEcrKT10970K9biS59swIBS+CulWHBkbZvAuU+iaNVOqN+q51IqpP
N6GL5CNQYi0rbMemypSsZJa91JrBjlu3AXNi8/pn+kSoCcBj/4bhBFu5IMFfJ+5g
UK3H6t66+v4X9QIBQsBXGhUjYF+HCsI+Rt+UKY966qHUDgb1jpnyOxZL1MG1EM5s
5UdIDoEwdg39xcoWvd8CEenLuCJ+aa5qyizF01SFHel+wH5R1F9olQEs32Zl+kJ2
S6LYAoqvPw4zXc9GobBsgAuQEL9xvYgo5pASDOKzlWXP7QnwAE7YY4eoroHWCMXk
ZmFncRCjcfD1ZqaQtIMM6KMILcxma0sdhLnJ4iWF5A4W5LZFawdzcKEX9arC+LvG
yXsaSj5VN32/lr3NsdgwIyJunBgObMKGi7V0j2JtrfRvsvr5wQ6bnYozGt1D+9Kp
Fh69zM1kbxMUTNxQv8D2Pg7XLDnqBkvLmFAK6srdoo0n04vtALsKhuZ1TxMmlypZ
d39VwdsKlgMXI2lZkjaX05tMucUU6ZmAK78DPTrmiNKZKYlYNSaJ3qRMkLqpDXlV
mYXluGk3UT0+VaeuCUoW+WMP8K36I+Yp24PtJmMic6aqcdrApoWOIOkr/Zo17jAx
XRhlgG3jJSpT/PLZrF15Y/18qDYBN3CniCF5q6baT3pfZU2VwcHE3QhnWIA+IXLi
PmVhHnbnrYz6bIrdx4xv/hb4xfH2eNCPKG8NF2zaslmUKFwExT9KQ7W16l+mBCe8
Mu8xvUghN3LdYEUK907Ni3Oxsdgjv3UlAKOZFJUrXIDm8GeqG/mWPD5fqYzmxe4l
PBgpe2T30MdMxr+PicnZuTQwbkjdlM/Ggz44afJzCZt2F9uNo5oMXg/MmCHejLlE
oIGUCPCfLrmUCq6apE+/vvzHU6zBgFQcuasHGfcoJjuqJXT5Fnq1jsw1+7uthnz6
/hW8mwUCZpnV1+9AW8lqldmNrntfV1wT5dlAIoBP5/eRX1a8ypWh6SrRtdC7InmW
MVrEvfE2QtV1IqxFeu+xhvhiva1bC81JF59Ttamf2LGJFcK60eJ9nA2c3nlOSgev
6pxx3wWaymeSqFxZ0sdfgLfKoFjsX98G8TyRFGrThrNvzE57BLs3KOYOezk7/61S
hoJBqmnPMvqPI4oqXx7hcZaBfryfwI5Wvvvrh1+Q+yaGwBwmLbTimiyJO5jgeJI5
xBKZGHRtDpCH4sxbN55AMwWtT18h8ZBODl3R6/Uvm6GYy751TTGELYAxFXgGigE0
Z0TBcyf5Iw3ZOKjy17FI04CoT7sOzh2xuGYP7k2dnfJZecBb6A+aFMC4QNGXhipq
/BYlNyOIm4vg2ixTlA+hvoaY+wKzAC1vOXARpcoXX1U171LlMbGhQYMx0UeK+i/1
f0Gwx8CApda91Qvr+95PK4OOAmGT+vJ4x8lgLHbwTEEDxNHNrXRQVBkSnndpQlmr
sxkvtD89vMwfG1RQtuEtvIQdeyA4rtZ8EmSTHl09vP6KEoufRRwBPVuxuzMbjwM4
hNjM8dRC41cy53Z7gRbYHy1y2hyrT7RKo8r2HPmdHvCxxaV1oFmpbc2AMOUpLyLc
cnT+aNhlxm+/pjPr1Drea0G9DvYAcBWhWSZlX+dBYdIdYZi78ovC7ugYN6cSOwMY
RGmZ/x321vwqkdddNy02UJ0hS4BzrPSv1nGPe/ZyaKu6FALCJBZSeXCNNxQKpIzM
s1LHk6yJ8v4bIii3htQzTQGXvG//HoeNgn4D9z6Cp5h4bv1Mac9XwuWmjEDpCgJ3
tJ5M25b862zOxbpHzFlO6RbYTuvkXvqa0/moudIQSnXBXOvcDmXE8ihIL05RNf0a
OIJsZL58Q9HfZkXa32qxTRME+ne9QDVE3ozA1gi7j5IeI916RLs1gRn122Xnt6kc
FRIxgbZ4uex3dNlxJIanMmlAbuxKHkw43xSH8DgkgpHoNMYIcuTL44AJR3H3YwCY
hLO2Hx6wx7akbrj6viS0O6dQBO1OVQNsY+BllwdHdeb9N9xs+mYJlY8UOWq0Msxi
abgN8VBbpn0mTA/GrlW35HrnCT2b0eqYzmPIav/+8uJYQvte9hMyr5sJ8+uyNUGD
dXOP5LBFpUqvA651mtiBdBzZVsr9Hg4ForGnsGCRwp14ANOIeTqpbLeCmEB6Nfr3
pWwOlmsriG+BlXWKN+62zh2LN+e8AHDFZTUGae9tDTwvnro06T6lYZR1Kfn7+6/p
UitDwm33N6jWkkppJdkXldGsLoBeYm9dg+TU6ciBv+0PEZO6bBenVZ7Czf5APYDw
B9nBY37l0FaJujHwE2KMg8apnHj4R0oHKBxvRAQV2nsV2FuyI6MP81RC7oUeUU1I
PiglpuA1xaA41VtCJ2FeErwyiHJQw7S9A4zODdY4yxeXrCn57+IW+yUR9zx7CLbn
Sa8oQy0uDyK1gCk0LpMD0rJ7Jgbz7cYayR8Icf+qsTcj8MMCQq0I3yln7du5fmTH
tkC9qC7QaK7jKugVJFukDwViEhxZNwLnZFcZfuUs44yhBkNuTHdYiOjyRpuMhtpL
rVMCRMwPDSjea6GRuAlmGqKgdn2ufm4veozxbKTPr+Ucy62sEV9SeCjpMJqjnEw6
mIZQNH/Fug/VNk5o4eK7XD7GFCwaSj+dvTa414zt3SvF/yUOP4YGIYczEqoUwK5h
akLotlK1ayL83KPQO0ZnqARMM5rP4BvOm5mhadQT7ed3oAOQHmeyEuhBP4N0xPtS
TDo2tr8E5+tiApPYuxj61nU1RCv1RX1zhcyFBN7BD8NE70TeChMVmkQECVACD2V/
rMdQyga/I4rIhekwl13tup5LRNXckzy3e5rV8ImwGiI9wqG16LPUgOfL80bQuIam
Vm2IsIPhQ8aZoloQtoaoc8Pf7CUPP7A6G5Oj0gu8nChOuzh8wJEG1VQGu9cZSSf0
kpeKW2jiOBStO1tgZJyPzjONy7oSLJ1L/dzz9PMRekg68k8II1XjBbxcI0tsSS5s
OJSxAbKTv76C+A5SHQaWs4HI3npahl7myw3KAAP6SZ5/i8eQETwAiU+AOEb5WKSn
C9rNdLguoBCqhJs7udrlSsDK7Rb+M79ShHyyt+ykU70c9IphkykPZD+fgTNj8/V8
ToqX4qmvKDpdU9gi7f4d2Lrm1Fs6GjBPxnBm/lbj6fK/IVBvV4fe9TkYsSFOZ0E2
cDpvkNhbVgfnKClsnaEJF7viKTP05MTEMxLDGYyWDPBQ5eVqBDbInWqL/5FNmC3M
uYUJZkTx8t2MbWxNKA6/7Qs8LduR5RuDm4rYM+48/q73gUoLU33UIK4/CF0yZXhg
6itptha5+Y9Fsq1r6UtmSvu17MHIn1q2+VSL9kv5ycsuRbW5CnHwKigqnhJhvL4x
KoJH6xt8EMMTJKi7n7yffe5Wa7RUV3Gw7thojr7PFsKR4QacRtUUigCNsOsBHulT
dguOzzuGYzq7YlSKINa+qC6Da1YK+XqXhJ6N3QMS1nqYJY1PhIOw6MPt+Yjl/jPU
NIIPaEO+gdluMn0YCKetMLUv9vrFvPoKvhidtaO6TlopqA41faeZWoN6IuBhKtb9
0WGPT62wW07JRIhEGo2SN1cGcOTqO8CQjHXj90BnlF9QQjXRddA+fJKPgLQplT8Y
8ZeHSEDpWKf4sKH3s3+zOH6epG4xnmFzC7bnikdJA/8uH2t7DqOwMfwGWOzSGxnX
pJnSjllp5X5fI2jutGTKYIg25uAUYweo1gO/zdKPHpZYHx5zphhAd5LvxM3OAxpl
zsRVGFwCNxZ/2cpkEbtTv/LQQTxQY3Nh9pChCSgocVf4ysz//7b/jP/kp62ucZAA
YnuyqPAw/GO/f4cR4I+sIltelY8x3klzb8H9o0/QLnQK+7Y5BgZ16wEq8O1y+5xp
vqEL68O7YwerZ7Fbj+dNdNpt4MaOPDExBYVAvOAu90kN0L8vjoY5WVJKBytNalJv
Ty8Hh9b7pHuOhv6gX5kmZ8edDGFbko6dcLAzLFpiEu9/IvF5Exs1VqUPAG+2d6Pt
E8h0jBmZ22YVFPNgh4+Ft3BbajLJAVwfrEsLSggSwqPUIeJ60P9MjvLoys3YZGdM
KMFJMIqEacdi1c48eem/Wb62fD+EDQOkKL1X9Rc1w+k5bkurnzTyE9t7K0TlVcfM
jrrdNpN1cXFnKdeHhZniLJU2zWLNdY+7rgPf1n6fyim1dEL0HEPbZA7vIuerNrW9
EMSQEGuBfbMhPdekfKcw21wEXjLFxLDA3hvwk2biSgRzmK22ZcIYZLgEH+UutFXh
YzPL/bGTNLlOm76rV2uzkt7sdb6kKSZG1Z4K80dAbcNwrr1MStgWMhQT4v0B4bM1
TZG8nh9QpjVW+hLJEJTBygqfijv1m+TjLHQtK5W+H3pTvo8T0rBMFF1A0Zm916Aa
cDN8fK85ukMmHOjmhvcCSXOs49hjKs4VrBeZeGnky6qWoi9h1IIeW0wqFMDKgRyh
zc1ps20Dy4Y05WbmHP4yZ2+U0QNUsJeVMu79o4PrjvCKQMfdICbB20WeaCn0uzCS
C+2zXJa/gBCSm39HA7IQHP31gv2PHA9lu3CWK7ONds2OMRdTYcWVSZD0eu+pi8KT
UDA5mRUb2PLBhKAjMX0TzNjy5KXJvzzXuuAlA/bDoZAnQ4iPScZ5aAT7OWxn2yQ2
0BA7iqAVOOb6I6aCRgVXTpvezOa3sRBMRwvGzOFDO2Trs7GaWSG62+8ke9AlW1k3
83JS2EF5xXPpt+0AeDuJ2atM6z0QGr+/v90AmQ8cirl5d/p0rge3ZrspaTnngJ3e
HxkYeyZ0PLy70/conC2QAOtUO0i32y+Ss4yRXoHQ7yqF78dAPqCtrV+0npruwvHs
TH9EIewkPiqNNuPZ6kfHgFBI6wDeMydIQpqduR9rA59Q74EKDxddNY6h7lbBqEQA
PwQxmYUzs18/7F9/Q6Ih1JpsoUe9eeMyihV4d1bu8kdkbkpWdJzElp1GwYqy9bvT
uBnRv2U+pPh2TRPRqDf36mTJdZGlkfdCj+mBKvzgG9M5EHP9PsRTrgWhV6j5jH5I
jdkZYH+mDAwQbbrm0q6pF65I1HZQvdZCNX9dtZgauKlmHZ3ioYDT+Bex/3rGB2pH
QbZ7Jwm8P3RLfihWvKhegJXEHc8YGim4pOuAl8/I2T2Wr/B94PSMf4dvLurPgfcz
SHF2Lnhk38jCbD3Ke1X6NQ4xxgHudhNg56/sJv48tVy+IZX8Z9ynPoFMmiQfZETp
5L96cd2X+U5kK7ZXbYiFBGpHenePr8MMkgpabfwiXeu4UM5P3iW9LTxnlAQnN8+H
LgcaVgKUrGsDJZElwgABj/ROqWRJSNru8HutiJ7DsAESC6n83RUhAgyPT2kyM357
kQHFZZ29g+jR1TWzkWsDAn60aDKvroHrVyYx5GRIYiKRS+/E+1Ccl9j7pfcAUQg9
HQvwmZQM0nGjuw1osISOLrcmfaYp1CXdNP6TYDnnU9mIONGCYOX7bQ3WuY71cgsL
4xHU/UYGw0MePGTdY354yu3geQI68PYyfziMt8zfQmJ70DKc3kTV/QVhjDcg5L2j
CqLuT2HUKv2ambcdUFip2XLI1RMrh02OvGhub2H1QDkVQugh+7leRWg9RlQsHAdx
lL0A1j4WFx1bw6dfE5yUvNJyaVwnKZXKHLrRUEGYAdxfoToyiCAs79eXm9ukFFpW
9r5yoYeabD09v6ZVSQkgEU97hpafqOVmK8TgaXy+TkXrp4TkCaWCEzm+k2iJvUA9
oAeEdW3DBvXfK+1aFVulsHu1xi6KccvzrKZMH5dYUvkL0oMKKVUYVIVWHIvgs4y5
LL301J5zQ9+tCkUd+mmlJRxtQCDk1tan/9HRgKR9nyB70Ug3vZnY5z2i6l3q/SQI
wspofljXPVPRnp2RkELF+0ay5579IdHFNgZcmz9HcOEcYwk6MdkKjRaL3kJNvAw1
zBBKBgHGIHletSp6YpDQ+fw2UFmKbPrUmNnGLB7dsH2WLfQ8MN5F6dkmXOFmH3m5
MC7ue5p/ZNnI4Ieodh2+9Zl07TEmFYQy3hJQ9o63dafs2U4bx+WNcwtjEgK3jsIl
suXaw8HNP2+q/urur9IGhLkEq/OA6ImHlFGCqNbXjIlCb/CvaVSdDS84x7kpFxjo
bOq4f4TTvLLyi0pCwzgRa6ug1ytbwOhnovR4zuoh16cIapMtBrA95VWsVVtao0W7
ekNdTCH7jNsIeCtV3RUcHwQAnvQhy+p/2FL19dpwMk8GajdY8LYjidrMkLxZnL1n
oN2S4bPhttH644v7hajndcM/GdCdKYTho3KEOpizyAXCeHf8GwUuGEHfDlkCWN6X
C787PC4pgA4fPLqHrnhoDZvRDIfEOBKV7hxtQb7Pcg/22p45DP/+xZr1oZlLvbFl
X9n6hJrmwuRoLfIT4An+gA5tHB/2nbec6X1++gkgtQGEFapdhMC0xsdhdyoAwNUM
uPLoDpg0lPUWpfFuKD+g9OdbGpmAVLc+TTh42LDjclXKCIfgXzBAQ0Ay+DvfoEKk
kOJUtf0WBEIxN8yKjhvhfz0ndUIFlGUpAVutdLiQ87ikvq72LxOtChN3rY9uJs6l
orVb768O58FmFuhdjwojkpQfuvVkpHXLjDsJNQ1XnjrvSvKNYjT/8I+slGfcawda
Y4Gi6gYSjQfEbPVWZVi+dXSnFctBfPw0NB0avKWUrwLcqNMqkQGhLiGyRjq4o2cA
bjC2YEO/T1jt1/MkUiHIz8ZTjnkqx54UQOcBtPJC+TdBlUx0AQZ7A5cRZuQmAp5/
ebusD9mmBHCjZuzOfUmhL/1timnq0Lth2tQkqgiJpc7h2sedTLpfU8UvTdz1LlSQ
o6KjYskw7HI4OhH0j/7B3dtu9+30BhUGWNOJ0ILocKpfNFD2ozfQ9eJdo8vN3WE7
WGtOz9KrfvpSXS3CjPHauwXcA61yGvoVVBvrjOELLX43gaPnBkZnp196IaoaYQSt
0KiV739KybwZ1EVPhFu+Ny2BY8XrE+8ca/OhpvajYvvi8bABGYYVQi4s3L4BR2+n
g6WRlkE23Too1k88+eouJzTKhNHTSHWHPdHfaUhHTEk44JcvkIdc18NyIqYG7QSR
+p9wWq4jnYgT3ewgpjK1VIUoNhPe7T7ectY/QCX/trh19NHoXJpgH1m+eio+ZZ4a
Y42FyNFHGStzb8Aia6Bmjyc7cmgPKLE3+4XJK2bDeJMMBjX9lMpaJhG1Tjq1yNpm
TXR74Tp9DWwbljf2L6i0AQVz+sMwZKkeFZwxQCnoB1H1zWRp0e7sTReltA5d9rdc
Ptj4dnY7xV0rH0Ik3+vQYgmvSeAGz7Qntsae8AyYI0eh5Vlz3dVnMs2rtdjnDwuA
tQQLf6X6FftgSxQXF9SSF9Z3tO8gffEhG7o5Ok4HaN1kZbN8K6CWUc4uSQgapCWZ
YwGun8eV9Fgd5bnk4YnAPwXz243eGBwdj27XeWQvOUtaM8wnc6J6wGTVzzWBZXGQ
LZiPiFDvl1BJ6CwdwCe4QFbDqiMUpGsi2gdO9b+x2i1kn96lJjco3wC4RuVUIueQ
atLdheDudy1JIxATLe+wLnsiVXUJ+LckMPpgj6A15LcD80ZdbITKMfrB1fGCiJ9U
bpqQsTNr+zxSrJlX0Zr0fTcfQOeEMRwTO/BsadXTPoWQEV4I4fD16GUZxcTJnuJm
SCxZQ2m6UAQvsUr0ok6I6QGuh8+IPF/zmzLPS20/80TgXZLDo7gpa+/OPwvBl/YJ
XcAQNyRCisT+qBzgBsLvjttHXXtWudxnPHP8UdQi2A2i2KzLVRrupKyP+4oSeDts
N4jRnKqBRiWSwFmc2UK0pxr1M1iLwqOo91XwZiFEGjDyFqg74AZNFp7t5gorydqH
qwUMj9S6H38XDFvRJn632Fsq3rhovfhuuvH4fDD3XI8BRPPXB4RdBgSVfWWSiLya
4PNcP6hiKQosNc48IW5GzEkDG0QD8J3OehMcIc+cB3KMk/jpLCkXaCygf9QhPfIy
YxZOI4yUiNeB+UoVgTCNy1FaKaA9NjHDrQhlxCzHSewOhGvplRQcHXujHJkianYZ
DZn1OL1MvRySsoFw14wWLa5d5sf+SHoxCi7EOCDoKYwXVJMwPsqCd8ZngE043sKb
qCraMYzT/GZL95NYc52DuE7XfuC/ojxwoPJzmHuGMDqqP6Mnja/FCF8Z5Zmbxm9h
wKss3+GcMWNRM4ONfJW49o34dIEnbTHMwOn4LHFBaPV+rBk26PEa7OyjaJoPeV/Z
BQpZuDGWIfwvxe6HEXPqSpLpZ4aB3tldZ4l8wnWJLPxEkBsz5WoK/ru9OPyXNgu0
vtkvgWT/vuDjmRnUGvngGop0omz3ioV2nbdx3VY1PRX1rXZ40NhAWb4qRB5m4GDF
pPoxy7AX/rxBSt/sghgutY3stOs/3sZBq1shDYZ24Ud1GWmYbHjmWOcJwRSWzIrA
YT3JPeBWhc2qu5+q3fEEuPSDwJCNFWJAdQ0cpMSH1OUpj7qkaM0o2RA5Kmnv4TiE
30SEW4uwa33YMnQj6br2qQTK2IWRXjRQftKzHO0PK4XEMcynqfMGxBfVUq7O6IGk
xrPYFtTiP1HC0/pmF0B+QjsbZNNuoBVh2QVzU2KsBAFws3c9qmW7m0s3irbeAG4A
W+hS9Mgf1J77EkeIkQhTfH+uilQYWAqnSGc6ReVOTi0+rvpm/lowBavY1iai+S4q
TKF+6tJqRH7k+vLPKqz6pi234t9IOEEz3KuNdRm4r6e7y2aEegmUtXE7sAGpk2td
Fzd0a8N0C7P8beQXMhgH09MmprT8x2EAC6vlvBt/qxpxYVvOKkzsLf1HfySWmZ5Z
Dx+QDbrNFtRaH/xDPa5Mjw89n1wMwxmQnV+z4lSIs0kk5Jp5VfZwRHMBmY9XvGL9
7O1vTWxXlm15uCRc0IHsKGI22pR11/E2364Bj1hhsIkpFvBInkdiP7d8y24/LnoT
/91ueefpXnWaY17Mnd1aSBYdXKRK+uUnnwxao2n3vYaONOstoZZL5x9A4a9Gh3pB
sNm6PVGtetigEOWI5kBvzzCpXfvPmdUXlGFek6r77BN8o+FSaTOK2fLDjInlDnzC
9IRcD3nftyEHtEQ59lIIRYDQ2p7fd3/pHiSW31wSRQsaSc23tXvJsLhdh3WkmGve
GGVvBt6snTrL+iPG20WT2A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TpJLGA/ZaL8I82xK2ypSYxIKk8lR7RranHr81FnQl9RKUdrVxGx6ZyzUIvC9SoBE
SOfx+3bdA5S9vwZ4rNEwGo1cuggjzLWsz/C9Y7i2OWIctNmlWJa4gt9AqrcCfKlZ
7ZQbjFzb5pFR5gsKkHJnxpkymBG+mliRoomFMvH0ufZQWv+AhUEz+cYOEYZHGvTq
GXqKd+0lAA9GhEX8ncJBkFLLn4SgnhTfDWM3J+drA5s/pb8w8S+DVyY94QiQKhrh
1LhgUbCc3HM6kMObOBRpZTQ75JxTvhlQBGXPBDUmVpi5+o/jqPCnB5MqE5/JTYf1
w4zjA8QU3SygtuoDQexzsA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3568 )
`pragma protect data_block
tbDUipGKixoj509nwcioIFJ7GL0te51DMvfU1x5SmRpgwoV7xVw88mUym9l3Wg+q
M3YwUFJui/brHBVqjHUAQKvbW/6baW2cQNYbSLdR356jfKm6ynWWFjrZvTkBIinJ
VV1/q8uxXzX3BsQW2PFFaFlsU3joOkc+KJDtVSQ9NIffh8yaQWAdk8D5VOnqpdNL
qq58aiIzU7MZ27Yu8Afr9wyMMHMyvD9CBcanxzt0VHGpzv2R5zYgT5Z7jdppD2U9
VXLjV8O/5UyHEf8b97m9wdXqrLrKK3V09tC+JIIvtKOTAPYTjXV60CNXk7cXIb0I
3CQg3nRePO6bqOIIM5PmnR4jSsJ2Tb6LtoydcURVGLGg5UFpIzQ7vp+QUcT9royj
IVJ6cJeG1H3R6biW6mOiMJN2payYZYzZrYVpKigSU5tGXec+K20LLNNnSse55Liq
qucKmqYVCWehN5TCwYc7Ajek9RXN3psMIP45bsEw4WI83i8L8eTXbEPvtDUWo2RS
/xgInBJiaJ16wlO9OkX88+kRxHxOVI9Ic01aR6t129tRnGQyOBaORMqNRjOOQpZ5
9st+bYgTtMeWhrUCRjKEKnrwcpDBYQMBbo7e/ms5v92gktnoKpB2hPJBFUZ2bB0h
6kKJlPk1fjiZBshwa8ECp5iT2ffQSH0R6G+3XIQffm9HpoxRVvslzr5aq2hc4AJv
4xSx+4MBNFgk4J3p5ZN32z0zukbwSRb1K5Qj7jtuD/vsOu/bmCTLWxkVdA9hXCVm
OIZamdkE9Zz6g+6mU34Ejf4pn/vdqkVLxt9LvHl96+J86Iv8pbWAHhuHqwpk5UuV
QUCGCFEVr1LTW4jTTmOTe1885pfqQdQw/JpymCjlZEO8x4TPc1LcomCre8AkZkLp
JA1SIoB8pCd5pLMVOZioCzGwoKu2b00iF6ErrmR/Xm6j6gK1xBvwV5asZK9p369A
spuOr1G0wOya+nfRtqrGTBbl+fcbrADTzCZuErhAh/u+Fr7ZxYKg6eLld+ZQ4s3U
QA0XynHu6/fS2BzCVvDbboMVzeHefm080jAe9xfFJ8X50BFNRDskCcJgQnVgIfdc
wAMYmZXtJDneAES6owgrW9AbZgSIeoe/Bs/d+7nbhMzhy57zsIEfV34+xyHhNVTA
kxDh35O+NR1CAzLrrOCIRL5UHfKp/i69Hi/GNZqSgl7YYfxTc6+lNypx1SFo5L2x
5frZDmDX5T4Lyx/x7dBTgJTnOa29C5TktF/3WMpqmPRide+TjgoymZ0kfDH9/lRv
4GduSWu4r9a8IKdYNONT1gqoXRwOrgSH6rXXWV4gTXEb1Uf9wA20u0Ojax4u/Z2t
SNSnSKJDxrUksb9eegr7REf3NWJTcMobbshNUZMCkohyElyqdxaZ6yWhWPQ4Eyck
+VYUw3OjzD3LRaj7Wtwv4IW+cJDAf7IoyYZbI4ET/qgz++IPa6yoGYvFQ8RXwxHq
FRWNdMyTIFfoD7DM9GcgT6mcM0i9/OE9zDaMRsolE4oq7JENKUAD1JGjdX/Y6s8p
0majWt4I56B/yXNc56XiVzEl23PipRY7dCCriCepczPUGC4JCtQ63zrcMSYe+8TV
LUBNMhYVMPs2nE1koqlRNU4VqX74DX/2SvAlYNRtA1DTwLZdldVtGfxysZvtkO/O
eawPEFk5rBN3yyMD1FRUqWDdmZGRC/306OpNTh1zu7jLLpxnZEND+adb/0s2zDeU
1YO4rLCmC5BYnUv8Sp6OsdBF3tdS8YL6+31773/utKRjwAHmZgDe2spOfcd4x5lV
7CvbIFMx0+2+d1Ssm0N5D++1fY5C3+lSMwTKeB9/IvS8BZy4CjGqBnNrGH9hdK+c
X+FdynRp6xnw/3ZAhra4F6RCbEEtKltNPtlGTvTxoRJV7sFj5tDC9hFlU1IFztiq
EDP17kyMg2Xoxy1JZbRgKBKNNIp0l9UDunPkP9+RDBUqIBHzJPgZo05LVOAv0Hwx
nEgY2sBkNt24pk2mj496eTCPUXcOyaQAqnw1tKYbozRHGRWP4dZjcXz+/6rXFzw3
V2Mpe47WebCE1YmxIom4vjc9yk1lmu9lNI5k9uBCmlo68wUUa6lzB3JbAqHfxZA8
op09iy87PtCDbHRT9cSCRTPmCHnY6v8OFpARFQLtEq3BNkIz1Hq6o+Sh7lmGB1hh
wQdwebJC5OsVVqyKU6hdiUnt0TTNaG3GAjSTaBOuRAWx5bC98iXA3t01uIdvw5Cu
7HQtCn4hfcqxY+lBG4bLLiE5VPJEwtM0Oftbwgv3N7UkurG7I9PYQabtNqq43tns
HhCmmHL62KI22cS1IdVod3oU2kjZwqsdwYMtUuTXxdrSUrTzdIVk8173ybQTY2dx
4/rRvN661gv6hCYOxCcZz51hPm8GqE4ZQFpXgg2O968tQ7Yk05sAgUjGV8gqXaDW
k1U2rM9svI8muVWyhUfF9IarmQ0ob4dNWQOmtYSOUIjpYmYhLhwaFxd8p8X7SyAp
b6x5V0okXmJSdQfBY2K6uOYJfS+bdcHVKfQ0oH1B4kRYiQjiit7z/IeNBDIoHsqb
jC+8SxUl5xl3niRSZXwBeBPMuWNSOTKej+lSrpbvhtfEmFhNK2kD3YZTQYE8lKvK
MjE+gTFfvnB4KrEiyd55eVWWIYiUgNdBZXLhvJ4VwC6UgoxLNl2hYa9brFVA20dq
U5f24+RGJ4kwbeQQT7FubpY4rjf+n4VGVpNDEylOkbFFDo9mTHrTMc4bYxKeKaM/
8x5ELI9mJIWAaurYTl8O8aAEim6r1jR7n91qv+6bJDWuvLMbqQColulsIzxrM19A
g2TNbMiPDbXfZNI4msjFUhWac8eVLuwyesa2/gLrfexYmG/z7ZX+pQyWhNROmuDI
XTJ2HUVPrhBVwQ6yCMcfRQeZGqCteYwQ8Tf/qfAPPjbRTAGCjaMlU7oE2WIyazJq
OQBMt9JZy5D6Z5Cy9Lr/J4DB9QiAlGo2TdpA+88F6UsLedDvr8F8eA/VHgx/hsUx
gFdvNn++DReeJ+QR9Ivh2PK3N0jLbHeJsCPaOUYJWWx2hfotnsVwHuTe7KrWVvNR
5UaD56XcEEeynooaCDhBvV6CpwK5VQ34ZGP+Lpft7P2nBkha6xtSuum7wa7EQIu/
aSAjh2rfeKoypfBdgv7hkl4eVxJYFKeybn96QrzMA5BlF21fSocyvljTjFuvhyAX
HiqGghPUE4K8g0Gxujjsese+G+THU8Z5MnAuqjoXVhr2ysIww64YmxkVu192Guh8
zICIk9r18qSFonFaxXgMBc5Z13GInvkk5YO2pWwEwkM6ANP2ii2iVcUYg4A7q1Xk
2Xpz/Y/dCGKKHe71hR4CwpG1FwDMvINEDnRATm6IoZ6aHno9i7WzA7VW1vXFgaZ+
3HqfU8BAJwm7PEshxGqtRbHS9FN9tfpnAoaoCzngOpIiyPgeoNpNecEzGESNzOC5
V1VzRYABFV6i00XzOUyJs1wsjP2mnqUHZ7UmSWxt/NV31BGQmzX3ERw68LomFUAg
+uIDbKpv1nrcROgFdtHnLuLIPIBs2fdIh61f5MpnstG4KdT+CgNNgdbV+1wWhqTZ
s9/BWFPaj0XddlVL4pnhWpkJrPludPKnG9dqMcZAsPdiJVaxOA5s2E5MSq3nLqAc
YIUfl78sYfQsM+Ip8T97KtbpQw2vzH24a/XkmsJNpda8gtrvSYoVLrsEjJmdVviD
H1wC2BAhcocrbaNRl4XjSTxSFhexvv8cMP8KwmUlJoL0HD/YY9GlbmfTLdlcV3PP
luog7mY4SVrIkp7oj88OGJVdZ42Gc98VDFGwk6W4B7RTlv3eofxiP9nEOU+JMubL
5Vm/2BZEUA8twp2tuSdPkDs6d+lFqGxwj4+IBshaNLf8ArbUq+7ipiEThojlNxpf
2EddGB+HXzOelP3wcsowjFOOoS721nUpjMFbs0iYPSB/fRwY3S/aDGR1oKf8SAjH
xfouMr5RGshKuqzERjx03X0bVrjUkJQg8QfAaX0GMWmH1eLVyQzR/TId/iI025VK
VL2wY0lgZ48sTghKpd7ZXojuR9ueHxmXejWw/3ugThdiaKozsbndglFpZfc2lGad
HKNNk5my/CtKlXgS0/BbUXawPXBLYV7Il3HLRPFtyYOG4H0Te/94YZlF17I04LpC
3P/iz4lwlbECF0I6nPz5EivbBkjSngPxsD4tRLaTRw4wR9gUthnX7QKbYBy/K5Fe
F6UengtLV8c9HfWontiPJ6io50VCE/Q5400lbSKhA/1rqT6wfaqmU3RRYbcLa3MW
etqPCOPNGlLX6JXYxxSdUM3Ga/X9zhygseVW7eAsnvfMv6x+Zjolid9JKUH4oeGB
XXJxkSigPTxwBRgdUnQeDBurficRdf1e+8vBoxdpXnjerER8TnQj2JvxrLaOc5Cg
qSG+VhyTVcqwochUaGJzAu5bp7BAnQVKUJG7W2QlWdsp5RpkBZaEkmCNc78pq6k2
IsXUg5fjyK9MEgCsun2jntMYEMiOWbG3qkiejyDZsKkzh6hl5ihnAVFsKR3kcUXr
E9nef/th/5Nxm20P9JFz6ug8O0qzqHqwohRjefoxnfrASTya83KlfZhj6XRwWgv1
DL4vJukV+HsdJW/xXCIKGdsVfj14nFXlKXxOYbkblsBTi6e3UjCJ2Wbcepc89JGi
xDUPkfLM+zJZ8d4lNVFpry7gL2bL4N7dVHhhsnzYaBgrb0TmUt7qis+Ozhwoq/np
p761BV/4HwAc4AUu8fE+Ng==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Dgr7vxZtKyENtrS3gw/hPfXMFVoMjZn8FrX/w+a9EnSXnL8uL5N33dRe0lDFxHlY
Os2IoIJgqU/hgCOK6Tic4/jZnCdFyEruMEiHJyZsPDzgZFnH8kSQgCx8MqEk9a0e
JBxwoFrUyhIMXZDFZRQP2DVZBBsGdHSynaWOn4lGaxnKLQzuJbgrPHaBbzy2StFm
jDLV8zpIapI9oT2JQDgV7/WluieBUTqvczVa2f6gEJyBJywEac5Is2ni2YOJ7CGY
V+FB6NdqwLk0OVlI8nzs6B9US0jP6WaxhF2NLkbAaQ04BD0aLGt+J4kiiU1vGjZl
MfFDnurAaKjN1qbWhBqnpg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 28624 )
`pragma protect data_block
m0M3Pisri9mhs87XoLzPMb4voB70OxU/SVwTo1zETGVwlECj+BJ17d/ByVGXqvYv
uRelCa9TIdhAfCOK9IO5FytQGhMBeJZDbIirsKHvWAV2SW2LahTSvj4w9K2UX9Cq
mPdemE3l5w1csjPXPgUPOuf3CuVq6AyUB0sCfbk7PXu+YG850Yl8sA/MMZ4VHlEU
D0d+CGAthBVK28ZMXlPEy7jAz90bewgVdBB0FRSl8112qKjGdz0GI/Pr/W7UBh1c
Lh1Fu3K+2upXQUByputRxUF13FCQUxRghX1S/iwRxdbp/bThpnzHBKBeEuQvkPP9
L7/YgSSqejWtfK339dvS4d/ATcfq/UoaEnI4k2/sdTDt0t+Zi5tGI69Ol1UZtjS4
QGGhU5e1UTle3vK8PQkN7JbqSJ7AgEwADQsi8ZnmncXbO8HyCVijz6DXYmIryAM1
CbWpmXXlxsZBZ1ubHkvW3RAPljdLE6Buv+d7K4APuEsnoGKjSIzLIv+bYiyQy24e
oQmdePp1NLOXb4VgicjlRNESA61SoRbfePvzUTGTdiw5d9E/V+TZS11rnzwOQL22
FxsrD4XPyGy1KC/zawOOZnniO76UPekeJZNNUz/pm8ZhpgS1d4/uIva9d3MT3kIB
pxqLJlzrln3g/0rDhzc5HefFVCmCRVRaWFDWMqFyjv6mKjI0hcKeDFFUpPociU6r
si9DyF/ozFhmd4EEXpKPWw6MRsrILBPAjJqufN15NMUrFYUvbYpETB7U4zcm920+
+5GvZgPFQl4355kljksSO7zR7Oi7fkIQCYkRu+PHmXHlgQyTtrbBoV6UgVMjIJKw
tTzLrR/TmB9Rj31MHkD+YAgKSFPWjS7z0uT+uHHKQ84ohX0cA2egtkzJyQWivDD2
vyY0LHvrnRBLjir+mwFFpi3y89NuqDMY1/OCAV+ht3kNbTAz3vg969iRsMwWtSje
vlTkesVd/ATvXP5g6UFmUkIaAQ2XE3r2xCKpDdcGef+x2OYzahO7Kv/mLJ0OA+xO
elCTyKWCXmsMtbPXg7xBcJiGjnMw1ANCtJawZE5I3KbbVittefcLEvvS53IjvhLV
lF1EwkuRgRmvHOWICrTPTdlBcLax5+RseED8vG45/kYVZZmYn0YU2rIu09SR4q/5
UUIjfVxF/0Qbh5MOFRRw04xDjbbseCKn9kwCxnNooMtxVdMTzjgMu64VCIoip4Mt
HioG1MiNZ760UZgWhMU6O4pvsLNiz11ino5czPHE5hona9whlf7D2+I7gTvZB4+N
XOTyUG9bwkeEBWFsJ8wgzkyMXc7ZdglVTe/+uZTLod/faFd6UaJOjdDWsbNIx75x
syGrbVYBCZBY+gTbDZG4zdo2AkQsL2OacbFYSJ4xygbbmsMyZ4yopMEitR9vHx11
0TqJmLNZ0hOmQvcY+yTOHpFRGahT8y2cxF5IpqLA4abjFcriDoPCETPQiZVS2IRE
AxBGzgk2+085eKgLm/o1reXDIcd0YMzo1tKDIx5j1JviwxuYXNEc0g2T7pMVdnrG
N1YTa4mzVWhvX3/kzCoKzuQ9pr/k9Ysl0yQXsQuP6R6FBRYoQQxZDibWR/1wGcJX
x7FG8muCGLPPQJ2dsOYYTe2j6JgH0jcsbvaXcoPC6m+VWaF5pghcq9n8ArZXSsjY
FCSBv6TQKTi6cwgcCxRleUp+FSAk6cnpd8Aol96afM3XfyNzXKTpWXCZD62U3Qpd
Dsmdvvd45F6ITNdvD6Tt5cCD777GhxBnGS9EUULPsK7PChOYBwLgXKOsHXkeK5pq
/brRnVSpUkT0M4gA71nIR8tw10mNokAoRVdq1iW66UXBM4TBaxhGSH1pU9E7op9b
FWuvhEhXYjPwX69Z4w7Jrt4vCrjybPR1aYJH4LBSvXzQ5+qPW+KwjmGkVyn2Hl3P
2B15hq2E0kcInLI8INj0lE7nSFOSSSQ51x9OH40o0IaiWHPxLvMLwkCydxGx+vul
PQwV3SzyYeOcOK9XfjZS63Gg2gfVbGJoVjGjWsqwWSUux4WmD3TkQPDeXhM8Oa0R
9vptBxmsrz+7ihEkD+ufUdGsBUyJiHH1xKwJJUeiY+qyD8aJ+jufAWBWEnESm1Dy
rn8bnxIKGwwp1dD+UYayhFKcqWV/4VZT+wletUqVKJtWi3gZtDumBIp5uAgXwIxW
rgA7MbBSWvjG85uUV6EIr5v5VovdumTIqz9IjA2TlmHF1Pu4ohsGYJ0QKcL2jZtC
MvQ8IjG3kwBlGPu/tSP7LO92AyxyZp8MSYkSGDbEhIoHpQM0973eIzqekp+BFQvz
hKM/PWatoFoTn+3HBGV+eDarJVjllpX8XCf4On8WRxWZIB5Xu3IvrV476Q2kT6FG
puP/vjI2rn3ObVfBVc4ZxZv3A3HW/PEC4ptAN+gBsNFUZsE4fNPas7iXNk9OTIDK
6GUWTN2YTsGugLJx9Jmuggegwavr8AlvWC+PLjFDe9BAKw8JtLXlyCx9xLMpGRAl
FCDFjRjC1UfhWwmq5L8okLhL02IbH2WhFifMnbuBCBF+dAcOwT9tVwxdlcsUocjk
TsbH9QM2fWsh1EwQPLbGp45yE0paYrQ3lZ5UseXGXwbpe+OXLYICgdnBZip0yV3d
JITq5pm05W2qWxb87TYcakI3xU+unwyZMSVbLPKIA4wUvSmV3I7T5sOc8O+vz1ew
QKTGBQJyT92PDFjsoXZIiT94CYXEt0YQ3FH9JE+FEoKLIK+4OQx+sTGHwkq+WbQ8
Ihd+/ANg1SsZCrczJ0HGAjfBWcNDOTdUaYCCAjM1Hz6AY8HO9J62m0F6SLL3ipEh
JN0Ptf9CoUK4sOlZJpJ1ZxXE8Q5Q6Np7eYFoiHUK0xT/leli2ejumYfH0Eq5G2r5
tk51NbWs5OTp3Jdsl+712I3aCv2fzALxoKqScCkySZE1iDGmWmzMxkJI5XhJnxWt
XVPg3BqsJ4JFnDZRW4dWwzxi8roZfW8BnAwe+XX/Dhi7JCNaIkPErfOuZDRA6ljo
MCswOPkfRCsZkgw74T6D6q2phNYO/uE9iCaij/RwE8NzMcsJ+bfECNeKIIWd1YZ3
E6DzoPBQdk7ShmjwTkw9YgtDUrdQD6yqcSVkoE/iU68pDxkpvyXuPhbGFxefW8CT
9kuR7o5bzEAr0uiywu9zbQ8f5+70oGMBazfW/mA7JSE/yGwNE5h6eiOq5mO0IwKE
oqx9PWVP6Y6HRXnLERA2GbFlV61yZ1KKXveWACWSJjNarx5i6mlZk6GetKhY5yht
Gu2gZLH3WnPfk+dqp4Uiobpe0tHyd8hIKjjkEJg3X4hlfcCa+RsMeiQT/SFSx0sV
AgKSUOudAz1swWc+GJmg+5cEOI1sXBkBxsTr+NlHkEFz/uLJdtrITKvnh8Di1Iw6
qkWLYw0+rkwMwx4CMITuU4d5XwNpFL+HSuMVmJjqXS/ynE8lITKiiAdVa7mSo5To
uPF5XCBAqoAApihp+59wFLFbjPWGPA9g+xoK4YkFSxHcYcEOungIOoN+pcGQ203F
hrXIu5gc3DFs7a7u23g/RhPt+q8j5QA17QqWlujFdDRXyV1Ut82X7kIl1EAFH7Uu
P7CLwXDQuSP+DDFDxpKQW7oRDdF891zj1ei4ZoRJnitP1Trz84StmBdLTuAGPDx+
JWJlTNDbuowq7F5G1Q81VWw1R3YbXzI/vIViOSMKv33OB6PIrv+9OYXbtV7pDM32
cNK7PRIgimcIq9X9szY21uNWd4J4QsvvZedPLgO9jLDaY8JTbZgBGa2y+3GyygWk
wEtDHjdJk6qWog180tqi79WosnSNTeGcrfrIrctiAXil2DyZisGfyCrlcjX1VA8L
AqYPuMrhSQjmbiy9UWK1bWt/ELWIMrD7A4TQI69Ea3/VgnPhLL4eUcTh06onOSW6
7tLuFf0U8hPEz/YN7ITjRp7KhPeXP5CWZbhNpkqJ6SSFhxdtrL4dE2Jr4irSidRd
l4gQnXmFREveAOwM+5SkSEe6L7ClVELeJhEcEtlh1nuM1xVV+GMXAwoHbm2vYoK4
BCEQWj+kES7UUnlPYhDO0mNacZugBbMzKSNHxnofbiImTYrLoUhYv4DJeSSRMzVw
IiWGr4kyJuig1Wjy1eLvrQslnxXHT30XnDRgEtY2qFY5viBtyqlQuQDTXJEe6AXp
orrBMG57Gf6fnvZtsCEFn0Od2OpYCRWY2Carl0Av+QTT0umMp24cq4au+qGKNdBo
WE9RnioQAnktZZ13rc0Vh36hFjmvARwFLKIzlss6hIsB25Bw4UH/AY6iKRnzfsVl
GX2rH39xb0crazdOxP5SQefYA6dFlpDNQFlWG6WX5OnrFdEdYfwjo0l6S6O2btxO
/aqiB1zOluLA+3ldfvjkEOXPHVxdFQl0oLqu12ua9TmPa/OaMz8xbEHn13AEYpQp
LbpfAiC/Krx71gII25jS/gLytBr18JTPQnZUO0OTAbtVKW4yGxJUoAfW7KdMz7ZS
vxmlTn8USHfcL1ziy8v/ru9QojvwkQ4jbW5m6oARP5wcax/lCeVdGDap4D8B2yew
J0uRJB2LYydKBN9+wkAbxGLrnIU3fjdKg644NvobLZdHftfEhnG2i9UabVyOTdfR
XGyuXpGjx3O3KoNvUV5OE0HGyM4APNvBu6ByxziZSP1jz2ZUnCrf11phK6GgV/0H
zAoQdZrMnoPYpPpQGXe4puEOxel023rcUsV4PaycrVHct85VsBppd0YngjQvxaIY
0fftSBqECLLVetgSJVEKkOfws/dsAjJg/AUAkwj+rxoBo6vbtJhXdSRTFiBsF98X
5HQV8DK9n6fVYTH7Or/hhuAsAf4s0X/gjcgazO2ChIPWiOHg9LnhPC6N6yLk4N7N
ITr+ERLRz0956+J79JOhxMJ+5RLfLVFJCCBp4K90//3TsYHP0ccy60AnqzsuSQCP
ocwUGDzZ627bSW/Rw/+AKaTpV1vl1cfzs8VKY11mS2eL4H3qsHY0Mzgtcvu3Z+jV
CqRF4+3yk9pPoG7QPansnDpJIjceLX7s23GsS2F5cZdcjaqQIKHBsqMKWq3iqVn1
ntUbv9hLHi8whaHQUHWjqD+kOiPDv08rVmvevu5FxnrpAE6pzrUpVz5aP51uwziH
8NC6K8xjlo8k0eYNyiN3StJm98jY88eLopIiyoFXcqpvMpZugeO3B6nc7jMglMOj
sPTSTUub6pcKzZextm+vxI4OqggH1kkqJgupHyQBfHWYFRHs5rMQMeojiVwIiJDA
HExMlOxkaJ/RoDtkMDrHPRcp3Rsu7tObl4xQTb8NjYGiWewBCM231WIDKRNc6VDn
PlrYS3D7syluSJhCfk59lsZ3OL5Avt7hSXBIF5TuknQsv60Di5qp9rf2U4CttGJ5
3GSQtQDMmt7l5UoFEquLDlZ6S5jwvLSboLyf6Xk8EhBok/M6sKW+DWPsh49ojFfc
t/m2ncloBsLPrsRg55xJgt5a22O6tgV0rTdFhcgZ0zPEqhgcYSwnwW8Oj/rjNero
uaCKNhtm+KxbBSt/EDGnLVLYohguj4bYdFvzPpkKXizoO1mEfWRwGF+Gsp2Jyn4k
v6sjGe5k/OX/4UPoyvmyMlr2VKybtHu5yyMqBSU3N1TKNukijTplsmUzrza7EQR4
Fz2AShuzkCFphcQvwVPCSY149L1wQGsEli0q/s3BcNC0BqEF8KT32fHcKvhavces
aX1inyxBAqVIodG07kPZplIqbpXX8T01M+/zL+NPfA6JJequGw03+u//DRrSxCgR
w0fzLjFo8LYg26QBmeNyKeG6y5I0QIeadt14PR/XZ3CsQiWV307sQNJfXzfLP5n8
XFQ9VZC6mPqYkaqb0KuRT/Tv72PhUWzh9sn8d1s0MPzs0tYOG3+ZSqaFlZ04A1+r
m/5Rd9U8Zhwmwe+yDFnIc8ORZQntS0/ngDSudK6z2+81mkcUziQpJ3nVj+4hpdhZ
TxDOqQW8xqWhvPr08QX9JPbaRjlsuspNvd7MTDamjA4KcNy+KiTt+mgElYHMZtMi
YrOfBiSH+byoXBjfMbopC985VBvTrfzfLMeokY9mT3BE4gfgs9ldWHSahg61PVWo
uJtmD5DS27duho8lKHbab/qtNAYqxss5B9BBPTy/BC9nxNlDEpI99px2kLZSPvAm
nF7Eari70yJdKJQQthP8lSHvjUaubhTorVJfUJBmhTn9KlOVCzE2ULBiGeSdUnol
IeF/dvwCzESH6fYOjbsf9LTlgKlp/Yz7Z2c5RhCtQrT1WtvgqULwT1m9tAocvbYm
p2QbPBlR/qb26mjz+LGBV8FuvGfnx1BaK/AUCEyCT+kKpNHFAXhYrWz0gy3BZhdO
l0XUEiYW2An4KQxGVFp+B16AcKlLBg+L7UvFNaERJgWlCRBga6a0d6ZjKv5cBDIe
wrRAHvV5bUZhI49ULfzE8qMlz9GblC9XbTnV6Xtt3x5sCmJ1LEl/+xLT5LxQEnSn
ePJtuXWPqXT8cOdwN7I/DDhiMXJQr+Ea9qgQ+cvNfLcdVGoGug2gloVaaI4JeBuj
qqiQrbM9K6qffLoCUZUiiZDpadHBpxPD2h9G74vhma2STfQw3JHJMZfC+cHC49Ml
bI78KmCFhU9DXz4axT8nt3E1hrJc6CZy0bwSJnSTgooi54O2S7Dn8bXXMlKqqATS
OvUsoICT7NQ7RwN+TXy0sKhvYB1CxLrsr4mnPPVP1gVoQBoX5+QHV1EOR8ITAc0o
ld/nTxSoaAoD+NbjnBEQVMnZ0ZqJWQFvspq3BOJjl9UmWIDGGKFPKWvBkcvgBJSt
UYO+fHyypxsU8Cq4QnCrCS1T7MI378kQaRFQPE/JY6K6IuEj5n0PYNleYVbvqUeB
8YvUUqYXPcVXNi6B50GzujG0Uq6q9U58z37FkMvv5coPE9wnZsTkpjmOjfwyuB9g
mZM2/liMuMTqEmYyZ5rAFCxqeCOo5i54p/ZNxDKjfbIIUcwmjT72hEFocCHkysVr
P8pZbanIr3B4opR9YjebhpAp+hFgN8wpXPR1ZRrber6/U/wkGbnNvxqcybb9Wcqr
OF+H3kpTVoVCGwSiCwhaWX6/CADCQiZFQk0x2q3+2sY4jnnBKrDfqPCszsFVr7VM
QEsXrOZBL53DobtxCx6qWDq3foSM6qc+DrGYerR7nZT0AEbKnNhzDrfKLchm6dag
zIsg/Qbu1dfhmqqtd9PPrXgNBrqqcsUAckcJ7R+fOoaIQRUP6fnaUEkfu4zh4Bfd
Xps4A/LBSzTiufXBqc272VDkjybpkl6pFacCuQ2BdkTYUvNqAZREYuZX3C1mVJFQ
AeufE60qFprt6RUSlZGw8tCxtInIUxPDWHN05YBv7PuCDsY59/EaYw0KBCsxw8cc
UIKCkIit9FWbCDpfflqh2pEBgkx3h+9JBr8bqqX8dJX/V8SV3ryTWJxmWibV7Akj
VXAAGoCJS9oxHEwfvW6jRiYp0D+sy5OiOO92a7dlUnw7dC6rto8krWf3G49lkt8e
DXB3kdAN87jgpTBEJukcX1F6Vq9m2JSLAAnKydsy3O3kg7CoLl56z7yWAp4m8KKB
utBSUKm608rPEuf7uVFnK3XtDPzHQsvN0TnMNLY6HXWt7assGfvtOtyxDLgzRLyx
wgiOB8GSEEF6/OV3mlf8cuu1HMCNcWU1roD42TJWfgAoMT9qjuyWyFpTccnr9Dq2
QE59YhTTCoQOrgaoVuh7nmJmjdpR0YoG8k/1y5U1KPo1EucdPjijdi0s9lMSkm6r
Z//Y7Y+zVjr4Sp1Xr9Pr5l7ir1lBXXQMVhTiJpupHQ5szLm72fRTHO/VUNZt00qq
SYLfdzg4mTdP10y+frM8E95MnAjtGQZnvquUICMKinpGDpBWLAEtO8obwK/NsvOs
jg+IcWJNubpZGyb5lqXYVNJl+DXgQL8/HjMIKOnt6k24JnaceCuRIjLFzI+ZiwQR
MPB4PltuECAb2UMUXTStfOtWINRLBl3woEZzgtkWQeN/bwkYYvPuLOtPIa3TD0Ty
SfQ0fx9X8g+87nMGyKuyiOQ7rIy+r18jszsevT0L/K9TmhYoQb55AwJJirfZgDhF
4vIouZunX2aQ2sLmlSHcCfAzZ8xCfg3QeDcvMnSoWaCDC66b27A8GZ77G9YMbmTO
Fg2RvdnHdMxOys1VqQc9aEvbtECF55xylm5ovRz1R3/HzshBL+MUK9fn2Zzo+GLF
1Dxu6T3Co7hkKS1oV1aOj6T0VxxIDfer1ah4+46K4Z+8PEWUJC4ZURaM0auMLcYd
zaeFNZIJ8+FdyHDi+Tn9QsxEM152SZwxdpeXd+SPV990Fcb8aTtjsvwJFLOfpd1H
vNdFzWoUd0oy6Yy/Y6fBwm/QC7UM22YOjVK4/9o2py0pDDwSMu6iAZzZ/NCLFAwT
/E5zcQr8ZYa0/Q7V6InyOauJzwJ7F6f2/eGp1kAtUZLt+CdCotrT+Lujxp2qtAli
1x/C5oMb3JepyKaMjOhxfMrOxk8QT9F3XaeERk359FNGDh5x7Vro7zvSzzJrVPh1
L/wXbBfMv4GONGe9i/SpS6qrCTvVg95KLwYDZjU6+0rAf9993LoTnEQRTxvhSanK
kQuPeTE3/tolndbEIETmCFzTp26UYp5z+04Ri47Cp1HZR+eW5GTyLvP1px54lfxn
brmhmptyqEfBW3kXV5kLOtZhCZu1evAEWp9XwUreZsvNJBZ6peYaG6/Nce2gnomM
BWGC58eH9xpbV7kbsj541UF6Qmd6bkv8QMHz58scMU2eJIWM3ugJ+m0jyEZcoPn0
nk/wZEjq1kC+Fk+vgcZee5MwJFAc+H2cbJqUhVrTMR+tBhhhB1d4+8pI0FSk8MOa
Qm74sVwPDey4ZLsWXCycivbUeaKOYDdFX/RCh3OwZ8opSzXewLXFgeiK+8gE0vnE
NvcR6I+W8mrsb97azGba0/6MZVOJ76cvOaY+CH5ZgUSErGaSW+wsMhLp8g/6Ely+
mmmvy5QKPOeEfSeAX5MnmtN1TZwyBLG96BxoMe9uh4DczIJuQipI803aiKZCEysK
HelqhuEb3ST6PY2je0qQG0XGA730FhE5Vmrit/YPQYugBxHXUEnhp13IntqW6nxO
Da82mVz7DecGEfJbD9a21UMjt8jFa5c8tEpttXC98dvcb7s9uy9cIPZSUt4InPOp
9ZE8cNrt2dZbhOAo+0Wepm04BLtDSG1CBKhl9VT/ClYRbj6JTbwRVHoLlDPXnL1A
92D/OZfyEVZUgjv384QOACQ6YELGSVfJovm5PzshfZdpTdMQfsC3dDTe71+h80Qz
UjyAkQA7nWC1VgykG/zW4ffEArityNHa36z+mbiNlt5zENaQREXMX7R7WFwc3jYO
sn4jjO7gA19PFlc4ILLfB53lwJmVRCkXm699RVa5z627GOdM8dQho1Bes+Fmf8I6
oXVjxVuYNj3BlvhnL9TlseoUkeiDu7sF/cNXm75LK1JvrCtbwCZaV9lqbKzyxXAG
VCtUzgY0unNEOm07CkSFiGWRia1/akfqbMs3FOTanmwY6xjWW1gwAG09ns3HX4ZK
r/cwwClddQBM17Ez0ZASgCIywRjswZ5Klhe35H7nbsQc/tEIPbCtSLAvA1PoB5ea
5lZdgiMWLSGu+xZDaNCdeRONL0WM2M5qUwni2vI3r4c96uFZD2pXkJx+Tb2b/Bj9
SdD4mMF+kN6r/J+MaA5B/PP0Z/U7UVsaOJyjrJT0jzLL6lFlK2ztoG0ciC5zoQLO
RrXOR+g6CppRDeFLsQROgAOBYUPdg514k5PhNbnbbY4WP7K+B6YJ0b1qHVYkG5ib
fwzCbcx5u54l5HPpo/kw8PHWdIrfeHbKtgtH2hwRaWE8i5IG9Up7CdSNIMMRVoHA
FN1qbPkSF0hYK0jM9I6qO57ckQKRXSTgCmBwud+BYcLpxkem6ZNPqz2q4ebLxIP/
X58Qqoay42UNF4mzNeqX8zbH6kXaWJReRhleAWpl0tzCT7XZktkoMUsFXKMNcT81
8p9TB724O1/14asH2d04UmKD0JAiiCjqVbMdMau4qWo/Iui4b9uBMUwYTBJVUSny
vWmNOcaAjjSOMxI8jchl3HIKnKMDcIS14e6HFVGnfz71GYfSw4mgkjlUCjbJCs2a
uteJfsQ0Riwcepqid4wZVcx6JZdTEQvNO0BCp+D9rj0QV4LckwvBv2UoHJYmFQC7
G2myPbOfjPoQo4mG5yizq2aP7kfh9C6yvQGZ705FDMvdMN1vBGKmBBdRCgFoAx2G
/4P48u6+CB6V9Y10eQo/TxjSsQdymidoj9O1rhcZzaLMIgjv14MXPjN69r3MZDV5
RLwoBz8udJV+LWfFiwArQ+JW/5SURrM6HosjGOZM3CTsnmeUzFXjY3BA6LqdVGt4
3XMaNfPhr1BNiNsLEfyFT413y8O2yyPmWgURGH3Lxs/IkY+NmZJN1YQCBX7/h31M
3JJMLRiMHbTBNBFnOcdCYKy2hJw0CHu3kN0++pF0UZBgeprp3IXdrv6hEm59Zvih
iG1BvpYtduKRSpD/zs5A8qhUtwmr5Ro8tzJOh1iM1us7VyERGt5/sbbjQTQd7AfW
UzhWkPHp6HzwIjz86AGPB89JTuTp4sNwAZsglGx2wnjXdElx5h7528LJ3TkmXTU1
s9o7TYmpvW0QmYi/3x8VMv7Vuoxm5FwaGoWj2Ko5XLkWTB2N2YC0XFRh6Ap5PlsP
SvJwQLdicje/php+Ouqlee62W5DUn5xcKl8tWfEKi0lLUs45crZGC6hzQ/gCVugA
matw0T+nazIVzkSOPTwQhmlk+stJmUCGUEgYOtnVIa3a1Vcl77mTokDIVEFHqfmo
O3+zY+pISjc7uDMFddOuzZaqRyFTjNc+fsHC1SUObbpJ/CDAnlOFkx7Ewk2gx8N0
5c82fvE2cIC6dTKGGFMadlcDATvpNzaifTatACjF0WyZA2Vz0+vMKKqMkg+CDdde
DEX/4QxHe/Gcj6dYXK+E2nI2h4CMx/YZn1gcC+YmGtX+ydGg92aa9uWfs3bCtHdt
gb2SyTMjWE7iDEUWwOW7vZvObVxGmMywywXgUl3LzWqRu+oF7tNqu6tUIE1wQd7L
T5o6cD+NhJV0wND8cpuEu094lZ2PoO/1J+unPdDxzQOLnJyvTj1dsfziCN+pgfCB
JKGf0wr2GWJxVZiN3kT4xI26NHJurjbRnYU+n6Bzvr7hfMeBXwq4dt0ge1HclAnr
LFzjK8X/gw3qgYsfBex0tTZiEXW50831LCX83YsPBisQQnHWFwbtTne/C6K7ALL0
byyi9TZqqQJIgEACuaeCPF7JgUYlREtIkN2AtU/Qv1dldB3OBWN7eTa3/HYbHCaA
UJMb9soqQktKErV2Zb3SgKA/eRsfT3XiGiqTnZUIMydatWE439VpCkxdl/ElQQR/
3lVzcpuDylBfsNeqAyKXRYuztVOjyJE7I0AgoAKryoKPzycuIrphlaIIeVNLWiIC
+tfoidjgWx4YHQGhcxlHTdqEoOYTi3JYDvGdun5N9aPJzwBSk4JNBpIbp4ju9rm8
F7xp0SBf3alSKCc8elfQapDTYWaPAhjnQEsA2Itep+bonjGh5Ugi8qPxWvQtfN6Q
kzzv2uydcpTXZDqgQqDNkB488u8mjMMRLlbzVMBt9GSRHrmqbC8fm5wekNFfWhHj
xVjIA0q1NsiZVJd2s6I6Lvaha1dEJVuzm1wbO2Fjv1Y8hpjz2EWAb+rlJ3jXx9PE
rn3KLz+rnvTjnr26aDsiDu1s47oFoB40gLj7aIfaqd9hsSQoA5cmw34/bAyfm/Uo
1bOR5+3k/okmrc8e5t7ewsRZzheIr81Jd6ZEYOyg5tdVFJUYIOgLwu737WPVlzdl
ahjYxq9NCAP0/7z7lJji6uo5ohYo5F4Vf5dIKIaE26m8Mq08FEyDzPjlro9EYqdf
va36R9FbKV9JQUHN8YPoZ6TwZHA3S8KU9TGkEj7UiHoWaaedzbLV2v2aWANWRpSh
PsY5q3KoMxBY0ZNPutaga98t2tnsW/SQFV3Zll/KwTAXj87HAk2XrxhZXx2tfYk/
XSkUwnHvoU4dKHZ74SbN207T8W+6nQKO2+EM1f4FQ09a0rFvfc+iEqR1yJFHLKOH
zJvouhbcu5ufXETnIxEehBXldRWF4NQMlNmP0/KrBeo1J8E42+4IqGi0uNLW9Fiy
5xc/JNb3PdyPFNOsLtn2UsRg5SpH8U0Ahdz6I4YRIt+ltT2q0sZ3y5Yvm0vA6mQ1
9eO37KdfCywoQxJtRk3pyMcKh8NN3DlUh4F05nkHdFrmCyPoGV4wTfyOxPKL0GYu
rieYQdjOOON7QsnU0v6PtMY8iBQBXWbMaFuLS/W3n38umpaXG2Fm2sgr9o2PNlw0
ObKVnTQuzI7YtWq91dbHaW5WoM+SZ8WJQt5tr1040s9DB0B0a6cwd1rqkVkc9iZZ
0nD7y8h7ZV1AKuekJb3owjJlrXnK+T6fU4tSypN/RtyeYxCAFlyDuBKEChnByHet
NpuDKhABcB0CJeem3SGpwGYvaAy3w+w2yRILy7wpG5AJVf1zhc3+ExukEmstb04J
mTB4+PZ8f4HWVFWnOaFNXA6VFmvpAbX26CfPsEOK/KvLSoUhJFr+MlHGtriaESK+
R7Y7ATuq5IeO6FSytMfPl3M0N/JaopZl1J+bf9o7zyC93LD9NXDEwQCY9X96xAT4
uSqK6jSlqIGufKzlOHBkDyb0x8u7vREfeNmQUG3sNVdHyzBwBQYVylXwvJ1pNDiz
7oxLEEz07H28Qn+ExNcQMOQCSRFVMGlyCmNhU+gCWMfdtXA1RPmVfIpPZ8UNqx1+
kEPHbJRaEcSRBWNxmP2wyo2S/tG79wmztxlFYz7T2cQGM3dQ8IOJFfrEy3m6IHa5
r0x1BuGGShmGrv/CA34YmpuEjfXHwMQ0aqffpSpTcOECQikpGyktHlUmlf5J8u5m
lj+2ROZRfxKm90iBE53qT7Mdwr3GJ/3VbdvCpiNzrsoW3A7Dr9wMjfvZUXnnpigI
VMfpfdLLdsBbFgulyZyyrmq1C0q3Gfe9b+isVPNtVzTB45lz4ajiFVqTO84UfjEn
iw9rVQSz03Nd/eRvt9eyFlw0j1t3ZMnutKQ6xdWRSuEextr5p7WEFYtVJg5NVzdt
G5f6RLnATdcmaBqrksoMom/YLyD41R9Y8/7v5vT+BviEof7F/kN04ht0XKzedmX3
QTLp4IVzE9Z6476mkRI/0Hft9V6t2nZI629h4ggQ3mxiaQuNvqvv5L8MX8eQxD+c
8iG0Y7HI4BSC+ScqcNmRYoUmz7dEJNHHGNuuVHmnBldbkgwiQvz2V6Ml1pJ59cH9
cBHtvECjLdHVvVcanaOcaoXMRDHoc2CZIIZcKZ+W63nvyb9B31pPNFDWujDVRvnJ
XB3sxTsMn/dNYbejQXxQzHg0BJd0RnBZErMV8c3p+GR85JE0zGGqk+jd5JYm2Bmk
2QCHTNbVDNnIS/ZLl7rQdFgLq3A2na6/4CzZbnvr7EaXVeATC9fnKjYjCMqWnJdn
VHhK5UClPWRaTpjj39Fx2b3e2+QAn11YQnOt3YjeWaNGCz7mDmI1SukuCGmUjPDO
jOlIbWneLoQCsZJPXdG2F0o8YBOrEwd4mRCqVgf28qADlY3pJRpSHkdIBTIO28on
Rkd54SQwPTBxvf+FjGpwdZecXggynitRXPUy/vC0x38Z7OBeTUned11gvEJo6Fkd
9etVXk+XfnxfIsoCBzynuYWmZGGlqMfp6Mae3/FAxQxXIVp19E37CYHF74saVuS2
o/G+ebKy7A7+qVTUBa/mXAJVVWzzKMfQgA7e47KX5gEWycmel19RVfa0jzrnbS+n
S8HzeEuZe3Mz2n29PGR6MIiOBd/Oid02p2C4jOal51XJpzi1BECUss/PXC1JA+i1
fQiF/i2Zocn96yNp1ln0AvmbsddyXxoXYO7wMV+K8OX1fOGOdltk4B5a91foSTcB
9zbv1qs2xWw0El5F2id7Lqm6/9l1/+p0tnVG4ViZL5TgWyQ8AAlnzLEMTisXRUtB
yCgqxtomYBHEYBDT8ZbPnAND9kOhb6xKS8cehlyNnK4VuFAkFGIFHVGAipTPstmz
mezgOHMlBqdR40fk2Pp7uaz9N1jtyS6SoICR7szPwCE8OTFefpDiIrU3/dEBnSOw
EqFfs31j6KRHXola7tbWFwZun66vvF6nP+GmxHl9xqlTKOBR79qMLpxN55nLXBQS
F+/1zgtk1zQtI8b44xih9h7nd35lDWxC0yPVQbGcwM4LgYsXdxU+37Kv1/d7wyGX
m3GtLry5Z7vw/r+oZrBCfu6M3GqgoBR4SZrdmxat+CvDlmFGrFdoJGQyOJNszF7a
iXciEeIy+vYxh1K8wddIYpqr25PXzClCWzZujCDgWVwUTk0zTpDqmdEcvfqbcoRf
aOl8mmcyDBKz4LYagViSaFBqUE86QnuDHyYLNufUi5GS/ed1zz1w+phiXEdrjdWK
WbJhegPmz5+A0uEj5wLj5/m/IF1bGAm4V+nCXfTpuP+72kmTsPQNxr64BOzYIflN
jfWJTmL/QAKNnPl50mlRsw3lD14WMbN3WWedoeeSXzRGKzAyaS/N9uhCJjaP9I0z
3Cr9ubAq8sF6Pr6RG90OmoAYVoGQCWXvt02TS/H7KuX3TGo7lfZncQEPUmABTItj
4VwP669KxK4g87pGswIaPDo/oG1b1bhEKKTZoBFq/FSBB+HEXhzlyhTNq6XcCqnT
DzJ1nwumIXzlXiB47DWJjveCxr8S0Bkhryq/yKOpkkDk9ASVQa1p1cnZ7RycaywL
8JeTw+ujjs/gC9SC9qqbTYfy5TlLvoh3xULN+PXg7/FiffmCgvb1xsq9dYdU9rBj
pCP72vNZkFYZIU1sSlD9J7CS+QiauWckj/I6gCzb+8nX9ynV5qzRrMOviaYjYET4
2y4kYBWq7mT7rK5u4O1UfXkDKJjFMljHtKnFNO0La33kg4kT+mak8t+TbrD1GYBo
LntpOgYr2mKydkWYW4AIdzDLs3fKPUDgXcMeSXV2O/teja/zyPsU6Ly6MrbLQchC
h0RAZJ7I7FItHkuo5QWzMYlYu1WDLS1gTXl4P5FfEGkT6dPrV2hT7SEjAS5JLI7t
9Np3fF6SENMncUlq0zEBcS4pzgJ7Vew9P69QBsrJgFCYWaSqupHwglg+bpm3qqco
nRQUc7R/NOhJrKbCpDIXkVYNQL2UiRv5hg7Cw62H1v/EzO6DnMtUqveuK4xwoafn
d6QIdrFj9CnRk+a2VWMhUwkyOIlhjpbaHNPHMOg/uFD+FRfj1kaVdQ+huxesimH4
wMKGmwSEx68k2bFIhI/QWq8DRTmDSAJTZKpb79x6BKJl6MHKDxmal0EyDL+3D8Q6
V5UxJaMNbCQXMSs6qAaESim/u8V/h9HbEg/zG+Z1puHlsmSoOSs6ymQGi3SJqZLx
noNe0n27lG/UTQh9sztr/HW6uK/2AuVgbYCgmRg+hwI2rrVAEoiAsqADYx60rRa+
95+PGx9fI/qi5Q4SvHRCavgpMM9aWTAtxWOuPYvJpMn13oZsVo//OOsK/rS3QGRV
M7YnQ1/jeKwdxkYrvEDtlziOMG91+IMma/mCLkhgP4d7CoLtlLHUOhsLbKpCJ41X
VxO9akQkUzIx0QNonLmSRlvM2jKLKz2/AnLOFfwsCEGFkzJPKiedtzFueTbhKgEC
EGIlKA2Tit8m+M3JM3B6avENLjbWlwWNQ0TGMgAgamuhs3q64kulgAOmL7oIcIfg
H5T5qRqtfHrW0Zb8Px28b+YpgRwr6+qZMECcIwPbi76jQX+dedgBV3Qao9GvFe00
MRbk90d+1tz4sMGh/KRsTBR6f668PxwaYqghz0W8zAlmZnTxuiXnzO7xeV3u49V+
HiI8m8Fp9IyjEbV/bLQi3EqYkDIFw0bvu0y74/VIKSV35f9XtTVJbYBClVoXy5dP
SgPSDhIIh++LzZttPUjcDaRE4lP9bsgJR52dOXKkpuRBUBw+2j1IK31kC1gh6Fd0
FXn33TJDw72WH3THU1n7UW+NEUNQNwp9YONklNIukd/XdAVD7n7GhfPDxvpFLEyC
UHFPpOrDYvDA+KahHAiJQEfkzlFPywj/kRBjs72v0SqciHJIFdpdAAlF3NDGt66z
XrfmoVcrnVSbXhpzNlWzOAmnDyOb7ZzdbheTyOp2TlvawA9AYJNGvSwnZYi4EU6r
L4lmrQLM7f8Tzlx6n8x6+qw7TmguAddeReEjlVv26V/qcEZEPe6ATMbD1UcxViAl
gNBzDb7peqHOWi3T8v5z2RrYC/SHInpO7/0emf4mdLNbF+ru2mhaECvF4TGjG3WI
zNEC27XJW9y01BpFE1167hTHKx6NtLaZFzh3KOMTvE8p3a84mOeADVrOaGbkCd09
vtoKdimXtmFVwgMcUAylkAlgFu1w/olzI+6IvKxVMMJXoW92mF0vM0sU/IAIFRsR
M4B9EuBYaDMB2jqu7ZB8D4j+j9dL7KxShfIe+RbyoKOlYQLi+J5YjeN18cG99q4n
8Fx4XaH/dnztH/gknETRfr8ts/ibp64kAp30tBmJl1qVT/Bk66cTNCohDvRA4tfr
HGPje1VRU7mcnfbXAf+eEwXXCqCG2LmpO+W+HaoaOwaTkbVlHvvESaGU3b8IUebL
+sna/PYWQTPLlnh8zf/M87EZd4IOL4uUiIZ2cjGdEWZPSNY4rtmjHRq9MREdF8u3
bVb83sjRA1UKrUQxtjH+co8/5AFGiDd7l9zBygQKDpnESrr10PmKjGYxSaL/Vphn
OWwnU/LDiQVTszPwFT6gvqoY94gsiOpUrlbcCETZyMClFypobkoge0fcVjrA0f1D
eRIgu44ELwaWk8sBhJUhoTHe85MlGQeqmDbUvopay+AzJ6skrl4B8mrzm60YqLHM
LDbELxHHm4jeGEsO/vKa2IQRCpD2bxRFgozYjjfMRf9Cff8CgB7exgKkoS2kTUTB
mINYU4cl5Rg2FZsH5liL0AMU5T8GUomuukVWOdtf8IUj/Po4Knz0ZH21pYg5ms0Y
cROfRSCsSdM8XawrJou1xmCVGVcCLY74Nsfx3HwWO96o30W6jm4Gl9ze04dOLe3h
xEx/yp+zOHjuH7qBEjfIwqqHb7cduRB3nFR0v/aH3DT028Djhd9a91l+SI9vLjUU
UGJEF8OL1FhVkYWJFPxmYkZwpWAdjS+b5XgxWStbXpT6ssHPCdb1kQnk9bXvOO1O
caKoW1HjlLw1gSTZQ71XtwwvItWzSpF48ZNokSyjF3NaWN5dYHacv/FA/gVbH2IU
ICAIP7zy8bYXlANrCnSpQx0QklWfQG3ZLtZuH9lPy2T3mmzE+zdavKaCswYaMkxJ
iq1Qhy4HLu0MmVD2zV5NkivcgRrOk1U7Nl+8B4m0mfcZKVHf/NZboSx8VUeCZ7BV
ddwvLxdQvXRlcDiVY3sg7V4Qbc3EOb2n5iNyysTN2enr4uHJYzjq3dKlJuY5YKGE
lyGWWZ8nuZ1V0TaRe2GWveHQmYrfv+ENfkqggJcsPCPaYu5vWZZv8UUwCE/sm6u2
DuNX/eaySGUd47rxEUJPuSFZuR2hvNDCf4ERpeSJY41HwA9SsdU7JUn3YHGbxd5H
xFJ6dBgljS8P4yCd2oZiXTcqJFiKOV5l+isrzsGI6/xmgOiQNo1neSvDniTSCzJt
6lnmXhV+6lIUMNRgMxr4ARX3SX3kRPwo7kGWhjjrfddovnZtG7i8Opn/DISL4Tjo
ZqR1PeLLY7dknVtj+pa/shbv/jNsX9LpszUMBZzX8gy3bUUDWkVhVshPUkHjmrM/
0rioh2BSgrnloCDXIuo9rUvn35HzUtGMJZCq2HTajB27jPEjlIhSjPuCEXgQGawG
LQdDyFZDYJ+VDojFMBdwZhNLUsT2o8xKwHNjz1LpB7sXoPBk74qDGAh6md8kn1Nt
8ctjoBmK3WxmKLFgM2fF9Lg6C+LRITZiCRkAo6FTG1OOG4QUY90Pm6bz+a/pbpjV
/ak6dBo1yltFeFi3sphIVeiVIhrMXdH4YbF3fo94ZQzO4z7qKnh+ITKcYWvDlBFp
ZHB3BVna6xl8EuQ+Yvhq01Pr4Q2FXOlo9ZvgAk4s58JEP5yKoOIqCQd4YRI2AuAC
vmrEF9la9AnIcm1Ow7pQajZKqGyksjiW+WaK5XdaEffXVxAmb3LiV5zpsfqAFKiM
VQ/o11VtTM4PpQGYV18sZpSgok7AsaRgbyzjWzjQRZqwQkcYKgrGYq8viiwICpN0
o+uqbZDuYkn6R1LPUi89e6yFuiZzp0sH+xfRsiFH09xDZP8mozv0Ax4HWphY6MzB
HWelfArMK0qfSwcIqJMbh/6zfLW9UGo9mC+8aQnh/GIO4MO7Ac9X8wdRwnCHYSRV
sGt0Ppa4cqGJ0GEjEddfEyzXL63+rCkul/S5F5hpGuGMSVZNfsYJo3SSooLvyjZ3
vovc6eZH/x4apXlc0rPfaOaONaa0A7E2r6RwTvhJnNOMh5D9mKPct7A7JiclhVbI
pk5hZSGO6raESw2+NmyyRnQs9Yyd7uszY0YrQkUoS7gBQzbyBMlNkdQUr3XZxdoM
vp5D1wBZC8kYnZ1NMrq+WHqhKWgcCQnvSBcF6DIpgZsrIwTsbCXab9xDawVssiwD
4Y0Slg1ycrCtpb3ekthoBKK4XQvsP6H/8KLJD7wMvsmainQ2xqXx5AIyvmZq1H/D
4oTHOwtqYDOQz4tN2mdE5bMU1za9QgLnU9vllNmooYx3LuESWb8CpUOP3EbNG4ix
Kk0CvAtNII9Eq9XawNtWYejcXmRSnwBwoIcSMpoyCRxolVFA+qqcxgTGMEOsn8+D
mtjEUqmCcPPxMG1gKGRVoDw/ykgWRAw8DkbkZXvrJscgZXVNB99Xq0rv8cTbAah5
FZ3l0waPTRc5f/FDgL1k94L/0d1u/Jt9SOkzsBX4Vklfpq1hsG34+MwfRsIBo0CL
Wsq0Nmg15i2rUsLyCnnrI5jA8ovtuh09xb6p09zVIYmvNyMq7LFOg9BiaAl6jcNq
HTIo8EJKchAsjms5PUlo+sNVOWu40pJSiCeT5vgm4yBb5CYY6kAAkwqnyaioxq1G
/DaEwX7Ish9UAQbV9AuUoSlYkzv7ERrmFe600281ANj9eA3C2A8XaHH87knY8CZb
HPvuAUjUUaJcZ2hy96Ig0PAS8e/gD0wYqFO3Jk28SksAkW7lKwPbIpQCdb9dJRLn
ZzCpGZxQwKfxVCCoGg4mm7l4XAUJOULKrVRE5VBXOVtruQKdPhbwIQE/d2nqZVQ6
llp+EPOhTZNcsksBUoqJv0QW5mlM42OQsqvbuWx4W6DXa/jMxClWNzNxmY8UoO0S
zFv2+NEwnpqYJa95PuDsH0GoSEHyueC0U0rt1WjKIIdJvQROJnpDif6sfLLGSRqL
tUF/r+QxFBHTXr8Gi7O2sghPyWkZ9ZUPANqeRkY7zzq7wJtAR97FVdZy/TNzAVYC
oP91KRf5Dql80l2szJ6qIGiOmEVAnRhJk9Z856zEUg+rGcywbCs+kf0iKnUlF5v4
k1oXn+/j6rTnODl1Jfhg35K43XGsFzQqExhszXxpobqLGdjBeUHV8tnPwn7tdEeo
1IDbEsW2/qUs/uCYxv0Zr+YEhhOxT+NxWzT/Jd/JyWcrfSo2difMuKaqWEE0/Ghn
lJvLiItzo246FgQwb7PUcaxsGqnque+iVN0AEpfu6jcEv4iacxjG62LyFF+lsPmj
DQ/yE83/tH6h32/+cDy56Xw8vNAdl52tYbomrao2jIlsLCY82bWoOWRXw7r+6F3Q
2ENiz1obt4eTKBnQ6fdCKI16Yxx7kL4VLkrm19v0GY1373wosDB3XKi0L+g+O4zn
lEHTj4eETRuDnzHL1aY6ayrb1H6MMa0EAKDXZ1EK+HKXQXmJvlWS+ymSkMt+m7ZH
rlrA8wEaPNU4iu+NvVaH9oY3BqPoqjxo58k68KikI80ogb2U7XjpViRhLyMTmq+G
+rLfMRJdU+n5f9R/QXrQWGtqqDo1DxlqLK53hTkk6l+v85I9+oY+pXZSBJFNhCPP
qo8Dhc1IcjzBDDyN2d8qpGEm2Egk7qpaOdeHsSBSuXMXsgH4dehE5m7cettt7/Nc
camsGJ8TrVx22Bt94eodKQqeCqU7nFuGW2CogvT7JIS/g6vfIv1wzgUNyIUjswdd
Ab4oDWE0gpiPhP0rdc8N1i6x9ihAimoHzJGAn4X2QebvEZqNKJ0nydnMkA/NfcpT
RYJrEujo6Izx8wa2v/4H0F1h1N0xukZRS4zhLW8Pm2OmgGQP1FpW3/0ETMqJlhC2
+xqNfTTfCwhYnoX866iQ5leyxyMvLMQi4EzPRLhanCmhJs/6eDHmbjxz7Ypu0qLC
EudBo4pMv2/+SlUHMjD9gcfgl7qyYuIEPfHFrc2EJ2K9Ggq23a5tKxVPQwYgp2m5
vd2beBulpp8LpUk1kCQejL4OrnqYeomVdo9umu1R9Dj+ec2mnCXQy7E8eioyu+pJ
0flbNEo/Xlry6s7mMFEPKrtj2YgD0o1Ao8awZOtqo7vJFhV2aC4rLu7kU6Bc+S2d
85O1cqUXHO6MO27siwOnYLSV4e74IQ5DY1jiIZn5bfpsQ4zaHpkn84t3YfoXiJ3T
53d2Mb6Osz7RHpyX9dEe5VVjLTpGCEt788WSmWrdP4uosPlcRENI/+5JvngsgL2v
WBnHiSTVUMZueJbi0ol08lbe/m+opwbpAYRzk5A477B1guUzU5297+LVQSK3U+Ii
vVYrruTgWW6oSLYW0HSlsYBXuGolX8INhwEMl3+Hv2T+fvihbl6zhdyHg0/9NlkC
wp1nCQ674uaXoTK8UwnmTwhcWSJARf3CiXfHYK5oo3zEcijeM8J51hU8sHHjDy7Y
0bzzd+m5p4ZXnR2PY9TEYKMgjU3oX/GMy4ml312cnEcvcMG6mvZ33z78Wg+RRZGE
8oLUp0KIvOcod7joHoK3Oh3sWI1i64Fqk4H0cV8kZ5Yb0e0Cvi8HDrTAhxze9q/k
smOx6snB9yWfq37sNqLIos2VbQSEiBkJWF/m/H6WdtobxMo8fuWlmXg5Ohw7E625
73ISnApOZNRvRZdk4ypZXMszyU8rajkt2uIi/YIiW8bjXRhBkH2VHi9DZXvupyzs
0q05hN6IgKOd+Wm7dmDH4qhf2i35JEPnRrQ19UhL0e731OcmTKq2OmrjIbM4MBNZ
POJNp9PkGNmdcjejpOVtt2CR9tg6LPMkM4MlG3S0JFEG1hGNzWMqvzIfG8xDHEMx
jrIOtjemljnlLqXyrrKjQdPHiriXP+AgzMXwbYYkMK6ecIdF4SrG0tVAet7uA1Yj
2nTSstIix4IH8G0YUWOLG5iJ1FK6PovBfamcbZqBtYTlpeVCA5JM8yYjDoDpIu9g
OHs6Jbs+7jxgnyYHW+6ZZJnfZNtehiDL6jEj8W/aKpy+XDOEsy/A0rVOeOLevLT3
gzpGtKoQIlMWTR54cx+6KWO2yTrAZgT/1CV+VOCICbL4ZKKCkxE7B3cRikXt5ah1
GaNWvkSC8a8d2r76EfMoIQCTFAF1GuUoOueSx4KDyg5mBrc1KgB1XOeUGZVMcNAp
rygRQKe57nWOcKfRnLsJtOEhBxF28ZXRbxbvzPHwxMEmlgfSJGtFRJ3zTiTOBjdG
lRfnmFhvTp50D7Yndwl0MDa2ObBA7bRVZEseZckMMWwcScBUji8Q27jPWc0gCZ02
Df17dbjN3GL2nBRM7L97s1cEZpOazuywnCK+3ExmLMCh15RW9fdxgnp99k8nmonQ
g1YenZFI1Yl0UbjwZSBlevjlknRKdyky+j/3l3KYSjTt1UCWljVCzzcuzWmoCk1y
IstX8h5y+pOT1EWzOSVwPP+M2pIeyL+R+ius+g2n0XBvosACf9EFmVxkjAxwvqXQ
pKVJMYemAkMhENAsRNlS0vJNfzlRcjO1LgGjoYd9CB/R2ulmaFbZVUPZIzZ/9+Mo
66cGb+zv/rRNcrvLw7jc88SSwDXqe2+ZLNeRxJhHQ507VgfnGUtxnuKNc6arz0tM
C/1PxlmbRVxQjOw+MtUk3yAQix/UyG2WWd7AR6uU3tZqYFBZG3KIEuyLnPG6XglS
Yf7J3Jn8p0WQi+AC1vN4Ajgy2WHgV/IyAVkfvgzb6wV8PDxKuWw5Hingde/14Ph2
IX7ePG/XqN572FNGeNAe4UEJkunvuIgCuUkOb17asQBj+3o3vteMDDYGXryS/nDJ
44wHFSd1XRvQs1i0cB+Tdz/0d00SyV4YB4kS9mNDlueSK20Z+kt8SGmjDQOoCePn
l9Z6OhcTNA4Ql6btZHPefFNazoIDHdtoDuKwBNltPObC89GPkkb5AgSYOpfHUFkO
IKOaZbYpKgSClzhdcRMWqVOhX1pP885ottI90BByoAdTp8YfHcJb03qpDA2CyFRi
Wu2TKHTefxolKvPbcppxoConK4nGdSPOkzoDtGMKhJdvcCfKf5wrd8UxAQvbs8Li
/rAXzhNIatmqiU2krvTN96yPqZPC96T64yfJBVv8GFseSmLupvmT+KelXzox245C
Ih9PvG+ITpoaZ/2Qnoh/LvqWf7FFf89Sa2PRaBu2yiihvYzYaUp5MdiP3WQe6t4d
sy4JZd4ZbYaU9Tr5PcZTD+XtdQ2NER/oi77XA5e0kkwhuUXD8ivl0sbD3yge17s1
rTOA1g69gQ8H0QX2UvvQy61dE4BLxF7xZ82Dh2sgyVVyTqB8V1/UwJVWK3aC/SE/
LaeMM9u8nkIk0+3b+Wq0uX7PM6W5Y4sv+zLIf6BHiWpvLfFRIMIW6tFg2mMwPibS
VVDtB+4LNKQZ5Sk113pEvAih5iHPtYZ5mLTINEWObNztabU88X8SOQqqEmfPYhcH
7vw0i+Ik2uHQh5oHpWYPSYqKVEl+EfIkLy+eQLYaSOisvs1SF3sg261GXbYDMqxZ
sd5mGm/mAq5GAmKNVtys2KvIZgSSk1xeH2Qv/dpfsh2cS6ZmCV1ssE9AVErwx+o2
0c/Mo3u7DuyEASQxjAJqPAdGlDkWEeGXnLitvDfEidqNZ9zO/xMgEWMB92mCp7j7
9USyzMDLfJfhABnZ+bnyMOwh2xKxFqL40YV/Kd9MeSZl4AOZqTXtwL4X8v9BPn6L
vprn8jYH+/YkkBoj9KQHefOXZsvELM8+W+CFirJ8Kg5oU5S4jlbw+NmvnerbEku1
K5+jSpKDXDAp8AVRZFCspSBbk1v/DZrd7YKij2X6kTIOmetUADUOVzGZCgAQF3eD
KAMxSKofv0uNSXF1eHscuYxSDmDdoiOwzYcfGZSOxIy73AyRo2zD+z3O/S0HnB/m
FEfo1ObaWkSDG5x7VGYMJnFdfP7WZThACKA5N8EziCuDMoix7Mc16ORw28IImjwI
rKsuUNiDfqwsFsk0yxu/7Hrg1dYIB2GpFlABauBJxjC28gIkxY2tC0/FyGt9xJDI
M7gcjcC/jT2RqVb2g3XDDZPfq7sw0g58T4rdt96+AxgCfE9iPY7Z1RVqueTNXWjg
jr6kEP0Do26lGK7yPdE9GGHmPHvi+wXVKsFTeamkkvyMA4XoLkBIFcu5oEBCtrib
F30JsbQitFl0pMclSmsjbH39dJhgZ3up3rSXtBgMH4lAxrCvrAIlEUol7Ylo51TM
yikPjyK4yxDrG5DRDJQZtljnEu/OVvVB0qDB9DQfTKZ7kZ7BeCTYkOcW2j3PY1JO
SWlFtGl5XFqlc9MaUy5ZWUARejEDNgBwwJzk8W01c05v4cngZcocCCaH/UVLaMNx
GDJ5/VxTpAk9FFenIq6Ct2abl7OHG02eLt91dNT/+OqCwTQ3hs8S16J/fWHNB8KV
mebpwcVmPD7pdBAiDl0//nPEsV/I0txd2VEUL8SX83kBdKbTdUwah6kYf92cYzdP
QiQWkb8S0IPCcIbMuRwNOCTpvo79AjQG30pudpE7rRzI353kK8xlPY1Lg+TfqSCf
F0va9tcavfI0xiRFuDEzeK41OtO/1WHOcKeh0/vjv+j5IKrzUwdSD5LW5voRYZbS
c5xLVDIZxnAPekNk8ZovufnrAkE6VrMC5q+3rPfAF+zWJLUqwQNCMHh7b/EBysk+
pr7vVAHvWoNLahlfYX+rnx1MuKtrw/R4u1iQLyAf6TwJBjgAhPvfpye7nd09yZgv
V1mKt6/mN5yPP5Ujnvu8Q4FGTvuqlxlyT+repO0EkM/t0/lwClRO3VBdAMtDSkkm
BVsG7tS4HiuyXggl8bel7RmxuTt9N4kKm6WBjNMavdJP8VUBymTKtMQBglai12F1
lQ5SB5uOOBH5ysxfDc5L00mvWjkGtsXQJ+ocITGAVSZtMjs1ZZXYehLOflodGzho
843+UgbFhOdbzQ7B0cKbCtDuTq5GgsdpmHb8chEZV9ejpuUTVE+CqEcRK91GBC0A
YTJlPVSyxNbVb0olcpDnS5OvtpMGhupiQDzJTcCK1HFV7vS07VbXY9akkp4FW18P
ro7Cu3MQtc8nlqetyuLlQMgf0h4eZJ6DsjrnvLTr0Vf+klvyEKO+ALdbRts/Dkq5
E8VnAAallU/340pbAQAtsMgWGiTkEF/+TTlYTsr/hqv5WImbZ8UDODJAlXmoN5NF
YQvanC3h7PF3zvSkRnYU+zlYOPYTR8b/DLFzIvKV7+G+fTE+l6H0k+y4FXZ1xrAe
Fae5/KEQFYXEQSbPYcMQ0nF3OfPibSyNOwMR+W8Swvb5f0zlrVGCCtFU6Lux4iV1
XKvjrwXLmMEi2X9ngD/Fd9DIHr71upTu7L5K3HOH5787BenjM26hsNrOdAo6nhZC
6HIyYtXVRcTrij83hSB6ZrV3YS0vOhf3m/3Yy0k9iyKzluuJ0s8ExwRHLjup9kAT
0nYEXrzoubqWp6g0GYRqlfsSD62Dy1hK6x2dXzvD9zu/PgFRPMwGGOrI0rwtkVvZ
Mo8fsRbizgOu/z7T90IFUbgdPz/GECugSV/krGKdHzp1B6pAsalGjPegiU0viYbH
5fOesn+PgEnW5+skv33FMb47poyLAbpg/AVZyVGto80TIwnuIn/nnIYug1Ggklc/
l4heucWWo+VFqjCXP87bvZEe21LxDbI2jT/Ja/FGxyozF0sOducK/mfbJyw3ZnHB
bOmHkjymImlYEzkn5mtKJsWUC1rB7vWZduolqDGZwnhY+c8lrIwAbrEdmStTSTRP
3Xgyl6koEG0s5LAsTscuDN8X3UH3Agf1AP0R7R6OwZ6No3errft/TMI1DC3I0IaH
fYeBAK1N0kBgJdFr1cMR0h8lhDC/Isdtr1dgp4JqMsNXk2v0MDI18ynmjnI97WV9
rn3uveTXimS9onraqKlcYTO3i63IKcHCGJtH5oBgVfQvprBrLtFY0R5GsgHrjZcJ
bORbJXme4t7OVH9xKyegs99LWMqSsj9VE9BOX06hN8mD4EwTOrPj5yXhkJtQoC71
+OAyn+OAMUwK/DtJjsq1+IOA9cR0Vn7StexFhHaHckpEbXvvYACwfaMRCVMC1CGO
DGlAtpuV+te5Xg/iPqIkyyZEayAWcsuUWqptBN7oxYxYZz6nerLoL3xhoyYEOcQ6
fq/tqFIiRT8nIxhXEEAaigzNuc3G9Xi/MjWw0+HrBFTx6b34j7Av0RsbazsuTOPR
vK/9SuDMTLbKkYFkthgeuAmrUnmemT42oTDZudqfDDcq3AGn0cmhxVM+FlhXdcqv
KsnYS0yEgoKXnhEqqOvG5sr3Pv3sQdZXCQEkDdNsSZNUxzrOJ5IXTLQvgyZ0ILKu
B1zvOJ5wmeg2C2S2fdYVDPx6eZ1nWEG6WfJ9nCxfXGIMRk/bnpCOPFcglIk9aKid
dNC4hBjqIdc9vIu29XoTSWyaesJHyhHT6rw94kUjH5PrP2hzOqPQwr0JvaOEEF4s
BlgNxf+wMETEzAO3mdLWZLcQhL1XHH5Cx9mm74PQreNgj+fRONLAV3doSCu6su95
nJti0OO0ZAu2SFggDyhzPAHcVn1YFcgPaswV/Mt1WGR+9JJrChbOEISHeRWwHfxJ
pjdIlZIXGk23dnj5N/4s9LRO472PtlJeoZWFOY9eRJaMjiPJjYRf4Yp7t65bWsuC
OVVvfxjjJcyYLq4ICZTPRagsSCZ/qNgwT8TUeoPqTeTMFBp4wUFkatgtAvHDmx9z
M3Cb3EccdbLWSDxWYP29c0hadRn7S/tLhtQ8MqMDbrFHHpw7eJtrMy7Edk23zCup
ROaIyU4cliNan8WsSoWDV06RjO4QP4dJd69K6xTkL6ehuCg+SFOLQ4hFAbooF1E8
hyqQtn58OdBL0rqOliFGO7IIEF9Bzx4djzjDjbruo+bjgeDcY30BjqX56WFH4MpJ
cBYR1+bXrBsEraMC/2tiY9JsK9brJZUJGBQQcp77vzgPoD1JYumPrM+oEKforJ7Q
asBbXAQ3IqL4aKNOHuMs+7eJkohbMHnLELJ73J/fxvrp2VowM/V/WN56j5RwQC3y
a0iwqH2zJ64HoGONdv/Wtw1pJLwxCs6Vrm1Y4EcgDbUF/S0VX/lYaj9IBD8lY6V6
mhx0N7TPflNctg8TpYD1mqor3qmLebjVXx1+XJzafRWvQ0zNX2xamSiIPJU2wQ9d
C5awGfO7qTXo4OuoXyulsqaMiMykpLHdrsl/BYXEqCv1KJrf3vj3kpSXZSM0SB7d
wLFoD4K3GRvnsRUlejMYrvxb1QvS944Q0Te9SabSj65/1I99cJNMqbknI6L8XX+i
qcbGy4GF3hISBiKOu7IbEbzxH2Hw23GH+q07HrQEsCSy1jRn2qHp+9O/FVxRPOV+
7g1JDDH6/Nsvuqq8vSwifi+TqCEqi/ANuqo36aTaso/BpT3MjoO+qKxwk6CrDAi0
wDW1WcZPUf1796sQhWhITT8Uzep4hwNO8jRmxq5dIEew3YJgxzu/p/fUQmOIjFVR
GqYhJarrrf8Q1hbHBB4ku3pqHQ4YmNN+kwwQMeLHW6FBCDJ8RRzmv7k34FdLMuIn
QidVSAfEmHllsmDCr9fv+pfLusbcl5loGOZaMhdaI5ew3Ks7uqF8SDRHb0rLtOPp
UjJoZl6DwSqoaNrU66PRy0ZXIL/8jzTBP2hlqQ00qlQzNyvW++joWURE1hflboZA
4D+K4RdjW9L7r+mQgJhhLeGXvHu+GVgIW/jrRc5tLoe9br/H99QsixAv02MPEA7Q
hWe+4c90YeAv/v83S7FXq9+08c5Uadx7NCymJISWm2w7HRPicQz9r8vM6vDg1PrJ
MiF0ogWYh6YM4EnNdYR+ewPcF4CEqZnG9S3F+vqnXTA6OwhtKj4DZuyB/7I/Ez+W
pjGKhIIge6sbwDUQk7IXvR7HlMSmBZ7p37J1GgDbsGYWXEpRjn/U1rp2Pv/y7IGf
5FAkucAvDXDZG9kFe0XG5+Xoa9BVVWwjkmahaQXvPjvgJSZS2Au3wBqR3npSGg+G
h46pvDKD+TuCvnNPUMg6GpGmFQAgMOMIigxcLoI5gJgbLc5k7Kh20KiWK7GgrYAl
zB2gvMOGPLdIB6G7PShT3nnXSZayliUO7QjJS4v97JWPBbvvecLQlSFTAbS/QqBZ
2MckDC22z+9lPYXG0bk5Aq0PzjW9i5zcRuKH4BytVdmUw89c73ep7sk+J0ZIRW5j
0Y6xNN9Q5pnvZsj1Ai4Xe0+OcOjlRtN8agBW0fDyMIXee0jCk9tgaoCEtswPJcXi
KXnb8qA2f5wUkMbJTuoopFVG2d9Eg7Xv9PS964f3Kytf3gy80cOGrrV05XV49+EK
qbPhX6sgvUEq3vXsGFfITbFvMlEBPqD3x2OxL50o8kvXnc1DECyFqM0KNhjiPbv8
4YU3NPnY7P3GZYFc3Z6hKRKlBOHlHqKO9op2TMvl4mfxc7bzbpAk6HjHybTtd5cH
zpE4dBxtrjON6JS+AZ392G9UZdfCZKqS0kxGX+kChkZAFgyW3YLnIRSbxg12sxCI
lqeC7vQWkbkXn5i8Ix1OjyL1SJnXbOOM+9Sosbpc2/n5Ft3Y0ZFlSviDrR5I7l5g
fVnJp5gHscYaj4j/ZNuD8Ba6+wYax52QwjrsJ662wJi884g5yWaOYHj65CGsmIWy
Vr24gr9E9APE7zrS8y2a84h9CibySP7J/SW2T18FXP4VI+mEQ3AQJF46mS9S2R6T
Im8VdqbAqiT/lqO0xfCKlgazXZw3TkI1mfwy9QH2XXw52xVl66Z5O8h1aPjsPhfP
5dA1sKPu1YrookY8VWAZCTUe1sZU0kwrhNfrBgA7bjQ3Ew11rnVX8S+5ttZ4W48B
8KuzPt9pGSRJJQkkC9UgtdbWeTyuUumhrGrvX0pzKa8P+CJcZUrQCS3ygkYTsT5B
xQTOs5HbR7od7xh5+TRLabbwa18VIgH+doaXmF6WsmxftRZhtgxzba26iINa/kab
Z2u/+yvut6DrI8GFbMfs2E/RJmmGDv9wNFyX11XmLM9r5+IwMAx+1jUntQcts4N5
e5u090ZYn17V4PpVIov53FQMA1TwAE5t63blhGXF26F5av6JMsWa/aoU0mo2jouD
bJ/RudPF5RZo7946/VyVCB+iETdJkKvs6K7dMC2rPsyA8LE+eSFxdhoms5R9Elt+
by8EwBdsyZmdzgFDnmUB2FXFk2athn75ze3FmstODX8FzW0d0KOckeUJmIqaDWPx
r/6YLGpca/esXDzk0Zl7Z0LemX32VPFEpfDNRYV4bqLuRW2YoNU16JLYZvJtPpf9
+obHKESLH77GdZzHHLmcFJP/QRldBg8Od5LGH8rYZ9VlnjJVj7I2evYgMSpt3+dM
iUb5fF62EBf3Q33tslp/hBEjt6RxAuuhIT3G9BmZMmVBq422vE/9VUZKQ3t1r00Y
0rtmNHpfJDFhsUTSG2q9DEyUOVqqJOngUwinA3FcEQ4X48EnouF0YecTeFiqc6/G
REsnyK0pmIOZGuRdA2eoF+HUIfW4COCb45GOvcKEvbUy6Smmzb6LBCyUgcCHA9aI
toAUhaB9A4FozEuZ9SCL6A+bhvUe45Je0jT/RJE0L2SW1l8LfYkMkn5BKWXaF9YC
4tNUD/SSuGMH0twO+22DqynHiLLphZjFqyAM2qPoDAEDca5ro6S7O/tNfdvAlPU4
WHk/YVTXfxwBdjI6Cfd8nwc55asBdBMHqpvTubreJfPN5K+4DaDZ9kROlFCkGyUd
hB6T4DcJDi8ITkJBE31OIZR13M8zSed35iYGAoPax+a8clNqupYl7IlF+efwx3hw
aRi7LkfWqlrP1ATzloRaqq66fBPQJzj7Gogds6t3wx3JKS3cAzXhO0ZuJPgvvtqZ
U28rGGmaUlk2vsMoRnEBLYi6HmNHUI4TSfmuu7ietOKTddP7I42xK+UoOof8/drO
zioFsprZvBX72/FQll1JdwWi0JfDmveVsrOdMX0jYL2A6GBY12yOkHNrmjZd+KCp
v+w8e1rKu4GmvGEBUGPuyofH2cRJ/I58gZMH5rmi2Yp6hX7MGINkawOA1lKJFx3R
yDoUNFAtLWMsLnfavd/WatSe/TlLU+AXM6/VpFC1a4qMt+5hrqPkgvL/szasJdoX
BzibzguLLqBmXKfXD5JYnC0oiG7CSp1HusA5HwFlO8WjDd55lde95xV4ddLVAOmZ
RlPTrGPtoAk82vuleHKiU4kpSd91FyMiQ+ilyIFuBkyKgdTdOhQUoQxCLvUgFh/j
Jy+PGEULJ27P/CYqoWp4eTgATKfPVJzVmEM+vbN5Y3daqVVcFm0qTInq9sFQgTK0
LO19tUd0GbgKgGTzAMDR3E4Dq933D+kbtMp8hkIPxYavUu3jlDLEl1KQ40u8Z1wG
okxZIiY0MsrKurLpHUQQ5dCn4yZBHRuQGvyrRgxrXxadthxau6t7V5rd8heBN9SX
IEmR5qKE/ygbvVFxffkY6t5WZD82SScSKQM8XPRDb+6KA4HVOm7SnnOdPGEpmG3T
h/Rqa1clDpCcGwHO7ealQSDz5OPLLxeZg07hnUT0dATISmCgTo9LiyvA4FVQl+Cb
AajrbkS+fsi5iMeeHRdf3bZJSN0VqrXkcKdDqs6c6GURvO+4X57KP4x7WzyLdHxo
g44Khv51vJ9VKq7Knlb8cd5vK8bsNqEX+f76v8UfOKrljRlKX9onApTZkAFckxxG
ir485OOkjCjVXskLCbyeOrPh78d/Ql7SqlZEWeolOcVPqtxwyQxMS50wgXDVXjBR
pMZ85CEUby4vtig9ORgSr9+F2QyQVZCubmRtUtwUuLfSm/gFItRu8MTR08UvK49P
Dqjx/MGizaatwR5Zt789sG9N61/r2zy0faTC+gjX+kMu1/LvB0J45/T/sKC2hYE0
p8VoWfeEqsl0rxXXW1+swsGL7WNN85bI+p8lF0Q2ffVekkxwJwp6OD06ifvNdb6O
i966uUxtEL/gdVWtz4v+Nj5xzhEX+oW10gX5lTIm1KgkOlYfshLpFKSqOfLOVzbR
XwvAKYMbx2bWNU4bPux91K8b/UQDF6Yfq12GGi9iS3YHGueL1twZd+J0+KScvK20
y4+rcsRDYBGFBLVg8F2h4mS+3hfm+gOVkLrvKDogck3wFD974FO3Y0/d5CnimxHe
V/pTYjMxJVnI1JiPQWC8O+Nqkzgv6ijMYYsPyRprdDpDL7CkQaqvq42Gnj6Tp4uB
/i5IsidyWaf1e+R63sxcRAkKqvIlQt3x8q56TwODA0ON891jPVlxpA3BQHUP/ef9
t6547Y+t194HfHshDnpjcxMfItvp0p9qZ9fjbQPVSTVUc5CNfNwNGKQOq73n0ZZl
C2TsMAf68ivvpb7fgbGbabhYUa3hjDH+bLU/s/xK/k/GuHrtonwS2/xCtM/VqxlD
KRyxHPWtjEGgZDdNXA5Hhdxtxd75I21ueU1JSUBZLVAPtIoGjKVEI+N6u957fMDd
6p45J4EdQW4hZvaTN9bW+kaVVnJ0JIcRrkUODiRs810tdtJlqmXz4VBxKPptm8CP
YWTm+RUpTsz8xRv3Smo/4XfeSLHcfWQCnk5+P54k+l/erXukJm/WkAsRLiGbjMqZ
EgOksH901iPWA7WI0A4SqU2oauyo7wQn9YBwh7+VUkWqoJ/MKS7l5o8NwqpxPF2H
BZKfizQJvzR/Dy5D9KsWDKOuD987NvBdSmxwJhJDnId0mtNoVAbVdudbdpGjoJ+v
/jrvrjRjrmpQ8afozIjamvNXLFAx0CWf8AFcNAr1faVPfcWZfRSSc6hgm8904qBf
vp/+3OJqd5Gk3ySZGQRzk6Fv6KJM8qejkz10RZRVlEb1tpSwARZq+RRlBZgF0AAc
9Omg7HKDN4inZHAHASQBspdRIrVI8rQb+h4NCJnzWXUQcjM4Rw0HrQ/L9tRE1f3I
2Xtav7wHRDaAdGkZ2oXZcAoO0Td+M2Xg80WtkhpE9iFo2yP5Q213WLjzlF2dwr22
bmqZcKuBLVJQNll1eGtIWqRJpZK1SjPx47suIZesBB2mSX8iP07PWJgvCA7yRoo8
26om7TfinzPdDSmupWH/SD6Cxo+0Pc3mSMAS1CSI+lGVYplMkFrXUvgOZLMR4aJv
pOsEVaybOfdQJFQdF7D8ie4BJb99sRLjiVLXZaSMcYpalVHiwrsmZKx4+UO8jWya
x3JPajNyMlynD/cv84/vV3mBLewJVhH3mAF3jCwSCtpETHOLPRjdaLfTZubeaiAs
qqUVxpPn0N4q+yHH/hhz5+BpCHmsL1iFTrb9EgzncvrfEgKTUvHfVnEKG9aMIrCw
ggk1rZsjvps+euKI6/y7nbRT/xbLiI4T7hNTw8xdUxy+5KiAQtJMpEE9H8ELMJJT
MUNwtQ5WkHHefcRC8WTpoXEVjdK3/3J5jXQSk5R8m9kFReXv8dVdXwzcRolNMabh
TLuIlyxIYpb/aU8UL9HOzO/DgH5ic1IZuPTf4L+sg8iHn8Hql+784BrCO2Se4Avh
RbctiEKeXeBITJkO0l3pb5QzQYZcsHPfxPm5VP8ao51iDTgxfP241WugnTdtfLP+
V4dcGhGpJdnwiasQgNOww+/WmhtKSXOeoMO2gA2fhbdLThL4/evYn+7xBjmuF4xb
zQMMjihPOA0QiQ/XPNT8ERSikDFC2JerNAldoUP8knh/tshuOX50Ii4L9z92m4Zn
POQ2BEDm+RuAvGDWCrB7lqWvYLmBhoLSZ9ouJkKUI2L4G9GWpAqFG+LCCz9unu+P
FGyIEPFwp9uFXqeONoZNF939iwuu77FI0GwnGLevIRPTO8uT4ODMp+Ks08mEYbiS
Owt2jsf/+6Df9Kc3edu1lCnvWDAJJ5OmTi76HX52jU09bjlkaKYN/J7VGJc5T/dm
DYd5p/zcWPahcZNn/Ns+Anvxp68PwuzeaXqC9brT9eYifuju7BrDFGHKxSKEHC9e
k7f71JePZQovOcbc64DS5SYTlPmYgZ1SBJM5l3MLKpZGtdOn7ELWWThcl8kcOx+N
rja9mbZnoafrvQkGAaY3/4URiCAKcETU1w/iqu5Pdz/x9QHYi/cQRKTd2PtPy9+/
CEVVsYZfTPqoAo9b+GU5SkLe4N+FVCP2KX3wwIy2EajlRnQ2DJCOV0l+4CgUYqGG
3eNItacOx0q0nEKrUr52nDJN2eFlZj5gFk+cQrAtDnGZ0jRySyWLxs9Ih3Mig+wi
jCFqf4+SMbv0AJjv6Zv89i5c1UBf7rg2VSawpDioNdn0uUBRFGvV4SSdjq4Zn0hG
zqcTfURnp/4HgWuUhwEzPQJs4E4dDBO0NUwL5t1CcdkWOMl10OvIV1Bl4d3a1E8A
plEVqmOHqpethW+2pi+G0bJdhkOiJfvmsN0FLCmUh81WbGgKfLu4jJ3Y5luM9mHz
f2NHVjzC84+g9WSK6dukbwAsqfq4ToRlXng6rCEMnMKIHwU5rt40PeWN9Ali9dBz
Jy4KIqAdAVFcDbDp1d/BSxuAMS07nq418ajhAzRxsGs2o0/EfQBsFwGOPpwfs6BC
gMS8S+nTPlix5Ea3/JDsDBJj6yn2rDxDtCY1rWdC+1s6HKyfReYjN5IdZI9oQx7A
VMhN6hQFi2OkeNjrEoA8VQB9mvYhz7APXHgZ4+Wm1+ZTtHRwwCxZoEV7WVGfU6bp
vy/DUh+Il3gHj70RQ2r0dxRPNJ7qUtaJwLuwDU6ecu6bDL6SuVJLVF3mmtwZ+P19
SxY5yvV3CIndntQc/laxid+1bLzR6kenFnsWV2VDqhmhB90oWFLwbgwDQFIhduY8
ZGWytV3pJiUlUu4QBaigkH4bg2Y48mC/guxFaBxQUGQeMM7+Et9p/ZW9dkvKVmVb
16BNkgdCP3uPxbUN7r9Za0qSv9wRR52GpupW6NX35qZfANVCW9tfbFltVY04VLuM
gC7Y+0h5MVfVa4rS/iT64VillfP1EFzXEcS5Rt8ZKgNpsdsG5+YYb6U/XbubL7g5
eRq2YK1NKwlJEJyXJM1LmZ4pnFe1R2TjgznaloupN0QpfVdmFhpBZWQOAyiKdC3n
28hul4BkjDCYRqwWgeWJHGMdlYKVgKRq4aUnUjJOMhkk4Kp6R25Xh7mefDoowu3R
6bQ8wA1hYbKIPTfcz+qSrCC2r9iSmtZ/Y2429zd4gu0DJbNzVSYkYVVLtm9qj64d
AIqn/+H6i1CAtrKGMTUkWpCCeij0nZLuFnxIsY2yiXHdadbKS4lLDqfCM2hFQU+F
3R6X84gS3ApE+mWyB1gQJlphmTyWG2xQdbbyHJhMk497o3ipeyiDPjSyCFXrAhSM
Vq0ZYmh/ln5nOhSNJFeniajWCJ43I3dFJHj1JIThPs4NeQwDMvjE6/Z0+hweBR89
8bOROVoeIoeFiRF4sg169o11gKuuFoIBT05i+BqzJ6R31QhbIjPQtxnCR5051m4c
AaDVbhb7smoHsy0ha3YAaSTtnB4f9hDQnQBXlwaOjPW8fqOmZqaqu77XGQKSWnNK
+oHuIXd4yzod8awd8k3J0E8XZhN2ISOXyeErgokiJgergDYdYoFfl+Y8mqxs9Pp6
sbmURicvkVVwZ1fb55evYlfXsI85vsVEDhNjxYJ6Ks7b1xMqYAsUxqUIsTE58Xz+
xFDMUQzEWQh2/xEi7juqWFmuaDCAKE4A4J+eTw54zoQPqgjcvTO1Moxc8eI6x8iL
9XGCyj0/MO3Uk3FoDRgdiaVPDgnYfp+fyWzb5/vYVawdb30Ej67P/4mhMIa9NGE/
sHV/NelGcTAf+zYQInxoFJDCzvX4TTDF9xG5daGozgwlCOmXbUNy0DVQXDdnZsay
545XzDq40Icgy04gsRiRNhS1LwCro5hk0WJHFNMSmKQwQUxCc60wavco+htVbjSD
k/5z/uqswq16eBPWBH+LwverjZnN8fQxZJZjd/h8Pi7XcUUSN/bLZAA+HUKtscNG
qaKTVYLlGGKPt2CHJ/CwXsFC/WMdeJdEQHdHCpc0adG5kMV3Pimn4TGh6B/BGRBh
NEaVhqE8kKN2kpCBwWve7rjndrfGJ1rnXfzvGrI1zTPj5IetjyGjPfrjRdnOznwh
jByKeKtilI+ipbd+x6LAZsrdgwKa9SHRYA6Bgrqrbgyv6c06iiTR9h9illabAJ4y
CptLnChaWDmLcM/L9sPX75fqfUtyCXlBf93AaRO04tJNwxhfoSoFn+FVVa4jXbv/
KaPcMnSE1sSpee+oSPEWQgUlO869EkNm8lW21dMlMMCfTwKQU2gzqXE2LTxndWaI
dHPAo/QIyuJZE596L/8NDxbUU0SCr5qdXh+YiiEnyMERFDCwwNkvIcN0HsHI5Ma4
A/62byjwTUjsdtUdl6NKfUZIlK/ylXgbvGwyyz6ToPEmQ3njx0vbrlMvSuIklEO3
uWUejq/LwuNE3OWPO5f4LGjE1h9qQcOgDXbIU5pXT6WxUR1oytej/zVtKJXUIbN8
YKqynsUJ4POuaDb+XfV9eKtnE0pifN7M1IP5366H/rrZXIvXe64yen3ydshhFvQ7
3UtjFXhREDUJAp4ezm6EcrljGN0+/kKkkEiUkGVh5rDEux+vHNjXfJ/8WSNZ444w
l6zR/zlvaZid/j5hBkEdjGXtsbVv5IR4GgUjm15wBpKLSi62DuV7skHJe/r4Q7g6
O0GTV01uoOMYS+G1AUTj65DvSt4jWziRm4SCTzRFafZpIekjQPF69GAicTAaqbiI
ajm5/CqLKHSjvS4UOIiTMT3hM+A/qITVzZbNes5Pb2uuDH3mely30e2DW2tG3JK2
HIOrlAq+Hfm/+r8O9nL1EH8COKhAdBm7qgge89j0utcUdN/du/pwfSbINKVviISB
jmi+WaEG6ZxEaGjfzgPKHwLii9W9VNn6bHZbZebRGGwBat0XXhbX7puCpnP2UfhI
ThG3TAtg+QrBuy/dwhJ12f3SyW5oqRmIHaNxgsyNu5YrTV3vLQB7KYr+FIkwkfVD
9FUChO2trNgKu58VXuYecKCRwxEjooMu2DgAejhqTx0PgENkiQEtf5bRKpJJPTk/
niCd5odd02ETGd/ORWqY41tQ0t8v0uiw89zNxXEgTiC+H16HeurUM8+BUE+9sjzl
8x3L9w/ZCbFFhfzd1n6PaNs96wjKLdI06grX94rHJgWRdwQaKPhWzfqwxSbC1Y9p
fdQ/6uB+Y6GELlmhzUaIxCtOH/3uR8ggsNmck5coZ2HUo4TJulgmCFw4hU/nC1Vv
3/p97apV2yX1Dv5sq3p93Byj1m/OY95w26gv13+crkG1NBs77E2HOAGIh8Ko0yO/
KiOWB79MjmQKHYwxRCy2OPHbVgb6hdyIeiTGmdYJPI+MuFlk//5eaWibd73WWSlP
ATNY+lKIs33704t8NME/3GxXfX4v3BaRDl1IknnXSiy9SMKuLzRwwwDhWABADZUR
PtPpDSev4Qtsxp/Q6Gi3GtmjmSNqaM9BIy5NWC+49GNpLPjKty8STLkG+kuECkCH
+007F4FZFzEEUXVlG1wZtSqx3u8UbTk2VefdYCrFyHcb4dpwiVNdMykIa0WozuXQ
eq8vlvdfWw+/YXiVZ/XvQ47k9LJ2E7wDGj73UpU0tUKru42WwmswBwxbC5dwNtxd
efjg3Wx/6GmXDD7W61iAw6wQc0jWlbBfiPwdbVOrlfVAAv9q0BOFjeITwi6TbIIz
hbEOOakGAiw9dKADRqmYWlSk1hfi44dhMmCoqJ+cP0dK59+TqYwVb3YRn33YTTkg
w6VpUne7rvk8Z+Rj9QYFnF6DDSc1ao7SQZiANv59zzn9PqKtFJgNJHdxo8MuewNC
1BFiD1NQ1hEGluQGJ1g9pcPmQMlCZppoI9DBo6T5WEtSKEApUKeu+679ZBBmz29D
vtTDGXYjdDYmckpRORWyleW8udosEHXTRSahj69iZyI31d2eXRiXY/rYM9A3tVjV
2jGgDioidVBb1mJCbEFk364NfNxFt5IIJnW28UtqmY+d9+vDCyQtRyj/55HXhfN9
QnsnVaKst+5BMgAaF1m9aLboA/pAemjmDsghSGnAW+V5Nznf1rYpW14Xuf5AD/h6
b2PffH+IX7vRv2X+ksJZYvKXgeMrwT6hJwvEvARj2jgSEQXUCAZEOgFzWuebnCQq
QmDwlnqhVor3d26se7OyBmx0eDmov3wg1+TAJc1295IYYIaFljxe5PAmnpDlcx+/
zqjSnA1uQ2e7A80pC6btvz1+ZblnrXorszyoF25GUyZTXkfAvQR4qh5O2huFOHCd
vKTBW+DqtFrm7GfxsEtlVO4LjPW4v5ZNLJ6B1Py3ELeeIvKlvbw9I8oxiAbqMYit
YKnXZP+Bl93rrrUioKY1mNatPlBWsEYuVhu6XE48+BXJcIa8ykaarSPUcS528BsY
bMYT8KZ+AzknUCUOlEdfhTMZV34aZKLA6NgsyECteq7q5X3FXVGpOpAAvnYXUmY4
3N3/mjzc6lizeFA/YkDmV/2GmUxWKNJEQLrhSPhite/ScPdEape5HrMeaNOqCG9Z
2nsbZjXYO/8wyu0qPX1ufNwSwY40Cq2otzJeKFyGe3xBYFyhaEqQAp19DNap7lWd
J1D2CoyvC/sQHa2OuHBH9Uq5KAMhsF9+VO6kcMkip9abgcBLpmojK7yDZrfZ7xX4
JRmPZUQuRt2sHg7GZ31rD/UBiD5BmkYRu2YeK7Dh/EOtM/4ckx1IpO7K2nn8YWD6
lkip6rvo1o3BaJBBmGydS8cXrQ//aCkPEOGtpd7ahPB7BIvdPKfSlJODHIcosTBA
gyZxNzzdNA7hCAz4hICwIlO5Uc1jLhklUivXmxyeYf1tOuh/qiTr+rmXl/r6Wmzw
w2TYKqR2YCpm1DtiloSfnbsBYK5aeZxQX7O6saKDiV9ax9wyHvBrRmfboD7cEV5+
/Cf0ktd/LoR84u/Yak5DHZMwg2C59gFg6PyftZ0ILNsJBamUc7KRIiM1/gc39jMB
1t7EDQE7vZtKykSP+huflH7T7x63hE/X+ZcVkdVQYmxY7lEznoFtOgZphGTJFQmH
HdgzJQVEQMNcAKXiWQ0jrRAwMt6F7cjOzbm3LLICF/TzYthhYwX4Uj/lnuEm47qF
njLLItn4y0sBKWk6WuAHQYnaJO4mqm45nCbTOu6fZAgz539dkdJVvlKu893vix03
11lnXWE4+kAnTcwgWFfomdnR1h5AOx1qHyT6iLLaoC4eUF3ry6RZPrFTh/oECYhC
2MKiivvEwTezy9UVnzJtOSXsdr1ANRiYZMk+HMAVnQQQNc8nMdvJ+aRwkWuHOpvV
EFKFvXAPvyGHo2/LRnIfipnwlkhAvKu/9OpGH0vd/EdXPkBHhNTaKhXQ+dxzM6y1
eKqymgP1F7rOZ9S/NB9m38brRdn57iBA0zY4DmpOwWxZPi7HcOxNZyKefDzF1Rrg
YLLP0Jt/OhUr79ClZzz6073FJg5CQ6pxNhJkW/KgGEKva1uzUzE//WgyktBetXpN
vHR9eokWmWX0sJSkTPnvKue779aC6xE2VWOGefhiiw0oQFk9KgpYWkLLhrMimheN
FijqNk2UbHKSvW/BRuhGzd05Cwr426vopzTvek7p7kTMTIsLe0JfNhN7kq+rWsiq
aPkQX52Y23dQ8Wyed1KaMfUQDcWnM7GvdbgpRJxhKy6NnCjCWP6mHmtBRpWRY40g
u5TyLo3Vi8y1Oc3iwNJ67OrM3xqQvwYz93yjRQYLXdp0oWlHUsGKa1XWi3lISVhG
eGNnCtdVdR+1D9wWzVD7sZhoEDswYTTtLnNM+Y3QSsOnvA633INAnxPpEDF+Voj5
+luybIWJ8RHtXkSm76ktUA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hHFDFizG1twVy4ScaGlvPnk0ELoEsGTZoVWhkq9rR1KY4frM9TeWfFwogh7irZAc
9WImhhd7GrCFn0m1ciziiisemLP6mIzraeMPehXPaxU3zdzPr9z3qZ821JMRk1Md
1qg0hhzTJrq45x20DQFqyLqdFZYKSrqdeDbIlwpaFsF9/hZVhch/SDlYp+i2arbH
YYXbOEu/G5nNl7PpL+2YjraCvgHIylEgD/EavjUZxLqNMofmnMbsIQNaiBtIaQVW
rZh3d2fzeSYiqR6sFf4VPF9xL1m7zG03lQm7uhuu0dS90xj6J3OPJ4R/WBdJp1yR
V6VcJBt8MT96CZOHxevW2g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 26016 )
`pragma protect data_block
7/X4BfzuXXsGRTwXrwzjJ5JdKXHXRmfwL/cH2yDEqrjy7mu8PjUqv94FGktnCLmx
nhlhK4RmInTeji5guq3NZ4JQdbYDf6yy6kwh6JH7WqhuSblNPAgGAie9eOtGnRtG
1W8O59Z3JzoFvGAgrOL6TOb8ih4PZvEpwOFvjxI2oRA9wlXyCdNXQT3zzOD07f3N
oMCSL3lITWgYzFNzdKGzFPkjliCrv1aOIUxsrZ4J92i+X41LNQ0g78GqKzQKTYz1
ktittTOfiIJX0FJaEw2edYQHKM70k7EKb3lw9samrVFjWceWB7hfm8V8BSHksp8P
XAfryeDXiFUQJtC9wSRwikizWZi8cWKzp7x2HdRY9CFDMtL/HDvIG5MBFDqmGD3t
S1gn+GXgKO8ugKVN+G0wFlfy0euHkXcU5q4lhVgXQmNth5fn7azmvtAOoapvpOqR
vfon2WLYL1Sux8pZd/9Dq0YsdZ/hn5nPag16zN9ubgJ9wvC7W0jLFhmo9ttIg5sJ
yaFRLQ75sMnxhePpC0j+60OMhlMYChvmBe8TvyTITPkn7YY7oqHQQAie+xnbHw3s
7gP4ttXt0oQb3vdhTYP0jzw9mrrLXWlxUFm2TR7OvJSsL24VijiZYe6JEUZdvoKR
7QEKZTgkTvLGh1xIC9aalROzUFRSishTcsItAlDR7S5GjYOcJJiQVwKKlG/CcL/a
LpfQsF7sul3m6DKgRMZYA9WBA5BbzsyGbuF5eCM+LcMvePUXEOiaKpUfbNnDsl4C
yWPcRd0mdGr3uGny5t34iOhYCxifneAavPnx9oQ2jBc7JcQ5PLG7CDMROKTcwg+T
cbUkaJuy3XRMOBOwwpA5SvNfVzkyL93HJNDFU8NQK6enHlIhuv6uWE2kWU6EUcV2
Jt9k5OQR/kVWvPLHJPMUyLsVYxV2r5Iy7P31Ba4cSb3NUAzHuGUazCKnpYj/xeC+
HhfCRatyWeITiXUDUlpLVBpcl/LJ43J8kj1XwK7l+GSLvuB+S5nlgmhsiwPdAOJQ
08umIQfQeD7xOYMYgTw0SggY439BhPxm6XeClBbK/w1jVd750htAX5a+E34p/gvk
GBSZ1n3i3/ASCq9OPkqPmUkcPiau3gXiU/04ePa47iUeP/0jEwLsNgnLj5FnwqFk
wZjmoiz7FuQyzsTWOh3L/ARBOSYBMJpnfHdJlYTTR4HIfaqRIZmSa9cJMUK3duPt
BsQ1yhML2AuNpVAiye60FPjOoNgDLc1TLSFmktdCkwNlSplhfzMvXmXzDrGtqaX1
P2MGmDKr5Ej5Eu8pzItvpi/VK+BEDi/JmuiNQ7TBKHPp/KjIEydztHkzuQE5RSKi
y74ZuyZjswe+r3ZGfOJjMnC/BpOUfqJGR5AAgImfDY0heAGtDirpRX17lq9a4OOg
HJHKp8E2o8uw6eTDdgMprzeicjhzyJKbG4jFh8hnSIIneuaFZmDTyxzfq1ck6Lk1
37+zzisIg3wz5JEmnlb0GjJLLRVFa7nH06Dt2dfAqG2REWekv3KGZc97jJ2FcTZI
zxpjI8U2sCqAKMThpcVPF2aLQQxBxMHGxZ1j9HJjAGtDrifAaDrdOaVXikJ+nVUY
eYkyMaAAex7DRp+539JobivxYI3QwRYG7Nznhai5E2cpJV6rb/KEazimOmimN57T
U/Tcnrfz6dQ+e7U/3GG1kIpRG9GG6oc6VEumIRP2g5dDLpuUu97jqnPhXZEVApuX
ynv6MV5nlM75Cq8V1w4ZEH3ph/HDmJI2LR+AI4ZzYawLaJfIlT2TZRIqPeew01Ed
C71p4UUjSQzzM4FfoDKheNn+I6VpVk5lDSrq82G/7gBXLDX1MAOMBms9ScUhrPSY
Yy5ceK7ubrwt6gKoGJq0GJJjlBmXPUcIlq8GA2inWNQdJmA3/ttRlA8hcJ8AYGCZ
v9Fy5JPDwElx8BEEGVyuolG4NtvHaTu16ewzSiYxOZVT0QI1Tku0dvt0TUqW0g8k
unW4G3KeAwsPpjDjqMMRxz603HtMiV6XRPUIvBJwKmmMTzXyFDDB3UdSlHUyQ4HX
u4gW5ztQCqii5G5wJBUXakYxbGNXC5DSDJQTDkAqV8i8JoCRaYl7wFGN256Q8XDB
o0wBxKfJMompdBYv+S/ySr0kcUeh6xnwM5vC4q4kfNBUT+7SC5cr14IaANDuwyPI
w7kFavReqAqPku5sUGtlVV3/K44i1LSFaCHDNo3ID6Mvo3s4fzopnkbtc+LFbgbO
pdO9nrQotPoDyn37z1IW4jc7i+BfmF6T8zxUE9mwyyqsKv9DHgi3X/QgUyISpO6r
nfxQRjhBI0M+sK3w+vyZLgYaCutBaOpLylbs4T1YeWs3DOPVsHplZpGVM9nzQ7i2
bwrCrKWv1LeQnTQYGV11sZ/HSXpVSsXkps5dHsgK3QnQM+lGhP4jppmkfE0TllK0
AwrLM7HDAi7hK47C2zfhFsJT8Q25FoWdJYoFfI3DaTDbPqFUElRpC+1pByvypJTJ
j2kFMk7YI9GGhEZ1Hp6jFeJqGD68NFR5LZBZ+5pyHRLt8d2s59zy1mZvxlD4WsVe
Yu21mZe5lUZ9IAcN7e7xXLyWXZL8zwuglPlZgUnrU5EAfesso3fm7EpRWPJ0FnZD
ESyF8vV+LEVC23QoXDZIjMPBHBwkbW0bOMYODXxO8BSUPKCLp0vl64MKSuKdm43T
DaKmPhcdZorwCqJnXEJaLdPh1VloNUfwEypPPoACSQV+x2QSsbZ5/m9uJff2QLDE
MJuOIBBvlXYwO/e/vg98EyMHsqnT0h2GVQPvxxkoMMqZo+Yezd3J6sAAzPGnV7xk
QTDQ81JkCdzO5n4ymqI6uraYcOs1XqzEkPgmBfIGsGBGYg38sQScUGPWl3EqE638
TNuG4J6PWR0Bnt2Kjx0SkZtIdhtPfWxD6hMbBC1fZ+zH/nrqWvdZ7EBOKHSGJsOU
LMS8jntRP0mMfIecFSU2yd7+SQ94S1lsj6B+BOf36qPfTK/UlaNM7mm1z6ylW8Ol
c1/SwTgnWmkWJdKPhXfaqwwgvJoT+wS0XHIf0S7IrIDTj5sH6SE2QcZbx9hASo+l
hoaVQEqkk6UL6p3TkT76UiGN6Xeu9iGDjS7zwHI22C2qjWhrIL1A9R7JqEWtQo17
sXggrZNp+oHUXqQkV8YOU90RtaDfST83EYbW4YsLjGDfRYZXdJ8QoJhBynw/MNGr
IvgksEh/NC3KSfvdAby9KOteIreYMEcC9/f6iJJ7vwdY4X11Jic95gqun1GqIgaM
+F9bQfRw0bRYbfgSUD4+LRVPO0gtunnhgJf312kP/OZLpO74/phisrAE8DnwfjFM
d9FLA2MHFrj5IsG3gGKRpIyV4NxDFisOgTh2jAzIORnqkLd1TDrPJXOC59s66bmH
IW5D43WYJQJpc/XoirbEb3JG/GjL0nNIFWEp/idI+lxPlL0LUgAurKF2ixVTNDLf
fxpikYci4rZWpbqnp8Pzrf9O/ioeZQeE0MfTnTsC8dDR9vIr2Bj1f9786HROQmMx
kameTIn/jYgt3aL4OA2nq+oDcLhrcnaMWqj+mT9/7++GlhcAF3ZguhjdkL6v3vh8
r6J208hi5s48ROL4APeCl8muWUWmb5+AOtQuUhZiy9vqTR8nxJpbajjPHS2Hmi04
6aosq+AZS/syxQlZJqWZ8cJYe5T+8Dx3+fzFIUL/tltN4Q/27OKUrEF+zz4GmiQ3
mUmoB7wWPF5hRVt8wq89HdqohupzUUQTd4Fhs4Kb+uvBG2iQTaqqGkMcrDTVZtkp
BIakM4wonL+XtGWOOs0YBO9QH+bncbGv1u/Oinxv6L/NHT29A8hDkQzBax+88686
C30SfnIS16NfSE3yeoaGzhMQI2aJvwb4S6/JFcweVwohJ0GNewHRVylH3+idnlBm
bCENpsDhOb+ajSk6PiQTkOObYF3BUZzRSf7JWmNLFDtk4aOzfhXXGTHpEu1du6ZB
4Lrw7iahQRwsQ1X2wc0xQ2jcysKkF0QrqpGRmZrFKrtW1iPI19fy4yVMrHfzCgXI
aN4ojngkRIE3GzN/7APqOYZcvrOOLA7QmVAWORxkzeE6dsXvg5k5atTQqUDThLXz
BOzsVNid9cwK+PyIF89/iAIaTOLsWD6/zhOTAt6oSfPtKZ3AOuDGd6TFGsf1RFp0
roAztZcT542y8XlBduJjc6byF6/uugxq18g2vGRyM/O7j39zQsKUCLMdzHNlg1Cv
/PWfZwe7aaykEl4qzxrDdqI/CRomKmLnPd/trBqcTvbVKVoxNp3DVsna2+yx/bm7
VG4Fg51nZiqMoKRgAqOspo+UZVNOTK8Qn92xJJkl8ixJ3QH/irM97iw6QsW+8Chy
DEpf5HL8WdlyvvqJz7H+TurH1OWqOqdSuh6dXF6ITEdx0ZznF4H8KxKGx4HnIdm1
iJZk8Rq1vyTkVg1WYz5mEVmtaKGK09jdz/JjWTwRACLEJdQvbdAp/df3ykUPMqIS
ybhLNuGcjjKDTZ9CZPHRGOpejCHG2EKNpKH2aW3v99QMwwqYvCVWzM+FsdahFGXM
qjTxmkiFJATvir2iqMNLdjEZtLdilJFktCnPh7LZZ7tkuF2unXKL7XG9bzk+TQa5
0XSRzvZLvSR+AASTHH8JJz7tSSFzzRd2TGYhmi4TQ5fhzPap1iRU1BePkST5T8uO
n2NBisHqNAASt3YzQde8G9Wfp2lu71YModH50obEVwxyJlWd0CfF79bHxDect5Wo
G/nZ7w3UhXxILD1wgL+0NT8eTAVORPvtgvFn/X+5+jhgKdduv0NguV0e3hrZ1ONZ
0TWEJ9OFtCW/zNIyVwbLe5ue+hzLvHgma3lBbpFJbxoRLHJolQFAek8l//wS6bwb
klaxX9/3IYXz+DM9BlGNs7DQqe+nEcXI7K5KdK0RWQwCT1mzse4UMV2t8PJPWaF0
AgY+xh/LL8DR0sh9K4ukEuZrTFz+ob5NmYFH2zhvWbpbgNLxqiyeUbLVmSRlhjfg
6ykx/bRLJfNLk0nNIqVumSh+tdo6f7vMuMiv4ixHW1SoOoe9/CdXHA+uxz315w2A
IMome16wP00t3SyS06B/ype7Yf/qz1cn6ZViBYOlf0qLm5WOgbZfQgU1jMKnagk6
EW+336VkxnAg92PT843rOduxmUk9RS/Y3llw3qMeMWlwihsI1Wr6gbOA9RULIozx
x0L1LiO1oLiDvBUX6MJLq8RyjhjKSfdcVTd+2ULTXtsDs1bjOGsy8B8pD+R8ZnJD
YiXlOB7COHbjJ9PJVoSbvksvv+NkYe1phZRpUfDdoN1csjoa0JnMyGUzmnW6BwoZ
zI4YdVR4MPLxc3GksjqHc8N5276ObeLGm2NYIQaai9t2Jo8lpFoYJ08bVanBN2os
xVLeQhL1yF0vbc/AekEeFzMKKkAlMbRuzI4MyuOX136l54X6ds/fFL4bd4ZqSDnI
EH7qmXsRHgfBtJ3sLy0soIRriAVtyTkxmlRgpg9NwYepHmnJrq5RSGAJQYu7CLzy
A3hhBBmCpFxkodELfWw30qoCtc97fbYxlzOdKbmT1K1ZVz3lY8TLydrmchz2Mq6N
+Qj/Q4i51ZwLcm+v7fkwq4UXqmnmJPV4P8atlhGPQWFf1O5GwIlWBB9EDVO52+C6
jBG5Ea5OX9yZAEr2E1sjaEUTtdpseHHJ796QaHgb+3YMzGKKJZaHegqiGHnh4kwb
fjvK8oDd8i2KB4LHZjeqEk60BIhOta9RlV0b22hQrqyW0qnXX2TSlRlCKq5LtWRe
5vMm0eKgbImhZ+2T5NgXuJq38ckk7bhMp4u28Ngod7yclnLVBfnSXnsvFZ8zYpNc
LALNzc6pJ8BWSITvBj1p+2MwOv8k9f7oxPGSrf4wpFk1JHDP+NoNvsA8RiNJR7rK
oPbev6vzwgZEr9DV9n63yFti+clXq7eqZVoGvI695AxSKYuchHie3UbrHZMZmYeS
irwhzEzNOzaqZ5R0tF5j8EquEqL/SKS/ZV4sqU0Kn7HYxuZVQV+bHYAqtJnrRoXv
t8FeTJVZRW1a8CjQbUSky/VMFNGG1NZzY3oyBUXVqSSrzce0HX997OF5Dkv7feVm
hDkSGWy84iWsYou+dUScpet8OnmHVFFPZBCmx3cfmeIXnSjvqfw9tl4AXBSQLI0/
w7psk7sJ4OjmDjO0NiQ8Ftgf5PnHVFR0BxwbUIfttiYZIcuFiszWQF+Gl2TCZSnc
+5IfPP9c68pz3XIN/rCz/0rmJ6TUKV0rLNPdbMFCYC6/ZQnCa2aBbucdOvhM62NN
ShWJYUKG2KEq4ds3dRfWcgH9Aw2gc2aocXNTJF/KmYlz/DB6MJ2CUEBMRfczr0zj
HDz6jbFcWm+pV4AI5K41KZgj9v6Qq7ItGi9OrcI0tZ2C5JwevQPvyy6zMP7iu8tg
5l+hKALGCLJn1Y5Fk9BvRFDBxQJRHOZMeg+fEE/k03hjLXpqCfOsZqTmH6Wykjde
xSkXubHyMU1ZtfkphaUmvnVF3m2H6MaYccElpuEi6ZMfar0SC5tqfGsrrCvRnHqe
fsP9PhmBAFCgQ0v6oNzYa41Vz0bsxpemGyilge0FjbzNwV61wNYlm6KymajdgZg/
8qe6YZdhzVvtdNB57rbLGj2E5b3wPwTZp9tzTg6/wo96N5a08iJkNwxatpV/VgER
yAPWnY1LdkI8JuOadjv13h0y7B2nqgOUGNi1vq/2zcIoEO0DuvpIXdll/cgcR285
dPnINXHjHbFrHlfFiLjGBRx+YgYUOXkfuTP9QdbHkJzbhY+M4l2mND0330vRgbHb
7CUWqkKIGY1hqUTx9gsVtoaERdSRt3DYvG5Ngoz7+pXQB2g5/k8yQRz/z3brEfoU
LiXV64AhOlK8KqjpbYXheeskdjnTCyEk3orlPf21GaODQdsX4DbSacN8Mq1y50Nm
xe5ogUxRUWR5BvCvYfslu0GLsTE7ve/pkcD3cZZpx6AVefsbqIxxIcg7jZlVI+fU
dsiPHJz2ScBr+uUc7hntbLqwXet5R93kjb1j4aV0L66Nm/rTLNnouIX7qhEtiRRx
9IZ6N+BYsZDOka/r68wBa0flJVk+MlOm1JvM7YNiBSVeUuyP5C3aUL+i2fJ9Cl1u
Trj5ofy9BtkmpzGV1yXHmJEPfKVbho3oPEpXSjL0WRxU/TQlTfi+uh4nIAgPLX7c
nMviul0mlW9Up7bmUXbuyC6KnOJyWo4QH6cyfN8Finp1HQFvutyFEtc3pJxqTnS9
yMW9kSOrdFYcWVwWnrRDihGvx1L/uM6M5EbA02KtTk8XCdgzYyhIgoBlmbrH2/3n
2Khc7R321/Yr+uUwtl2fe4LisczvEXBgM8lx/HnJMgpLNadIWuRrPwiL+OVVkYpw
kmpOBt60ZlWo9HEOPfBkzGkBXHmmOmFnJZ8wjDcTPadKK+6NwQB06FFSZ+yi91he
s+IxEo6+h+Yr/watgwyHBJ8PwY2Ox/Fuuhk9XQOzMVhuLTxsfZhfuj4/ob2gbMVa
gTuYSqoXbSfkL2+NOGlwuyKlBhqvnXsg/N/R2Z45F1urXrF5P6JayoQVAooGknx1
aXA9+8upR/5dEZV0Oc+LoD2gx4kcMgOFVc8wX/dhgtKtKSuleD07BfH3MkzT6imT
bUqD5OoUZjQMS9/9i3XOqlf8VH69Lrcw4BSzYO3Er7VRSVnGsMtbus+5r+Bd+4rX
70VIi84X2So9MUX3FKyH/zVfkyEmMs2A8prRAF5GD+n7p+xI3g9rZUFlH1HaBrdR
hCpvxQK1QZcc2WCJJ1FzSU/0crol+MV1zMP3y4mus5JKhk0tZcv5Qum9fQUZK2Ji
A2Vh7dqrzMHpYWF08nbL/MgiYUC36f6xQSy512gS0wInGLnqdld9u+ZnazLg80F6
XUPUaggycjVPTCr9fiK02N24GMzqCCvBl7fO0xMWBvTfGlWW3KxOcEAu3PRVe6dt
NcpCoxOg4wuxkxZMwP8+nxr39PD1KR9EN527hTmwZy5V2RfITaBP/vWARgFhaw/+
TGNwAQXi04fEcjnhoaFaOdDhZ0NYR3b+sEbpDEu6cK/ecXSemPSbuFGHS4l+NiDa
XG+2buW4x+H1JhuX7WvwAUNmuqMvFTWyymCS8Q9Q6/shBbKp4STroXuuj9Pf+5kk
qx3/5x0cJUblModxiDV9aUJR9i44bxO1Gvk5PWjLuR5eyJ8yNeE/CxmUEdpsWSbD
zkhKuBwELlVDF/tGft1DciQ8H3lz56315y9hcCHo7TJXbqsNP+Czp6Xygvi+DxYT
Ix849o0QPvyxD5w8eYMdWNxY49dC28ARrLjywN1z60bpvO4Xg0U05+CvW5gGp/PI
C1iAthDfJ2XmhsggW/5LJt9D43aG6SiZl8Fztb+ZrWL3uTMoe+y+zdEtkBKSYAR8
1n/sxEjT3VNIWvEYxn7UrA5HtXWe550JVSLnCgrm9u/nR/5BHgJPXZG/ppxtVx5o
vtVkY2Kl6iAFACaXqQ/KjQhun1UPKjHkHBqZOIE7HPiSfx3kbo/IlCkasq3Qepas
d4GqCtJjx1gHKNy8X59iDL3RAiDJQ8pXJRMBrjSCVudbpvtFMnkqPFs25ZZniNj4
RbbXwIDgoFhGtU1kP1vxGbtUvg9WTVEm3xWFF2oCNlepnPwxRc82zWFV/O4J4VyO
q0YC9vNaMu8rnG6icCALOmW56Pu6KEdN/cOniMerLSMwgRE+bDosSel2AQqBuvCw
cVI+2jRY3MTVLSJWx8kT4IaTJsFLL1SvY5g52iuChjH/ckkZAVOupBoe3qMmRGYK
oZtJp+3aTIOj2If0Np/++ma7R33my+AdSQGXPKerxGW3A1BOBatmyGxZlcVfkFC4
D8dPVdPSmweiUyz5zd46rLsWIdSiqokepqvmkpVb2oOdF+9qtS9AA/n1BrT7+6SR
6YUNPfuHkqZ/qgeyd5qzwjI0hOxCYRsmNhTzEqvJSvfExRmZ4WeBIcPULMwT+fyK
g7cOIFSwj2/gfFvUEn8+HZDaAM2sI+7OG3qtR2QaGdi+V4h6tUhcDfVCAVK1G7Rc
MJ/3wNOqyzQB0pHBdmgMkiS4fQThvfDjEsoGaCDmruI2/LRXR0pQoZXebUgluorE
WawEhrMpOzJhH+UoLRDYSMEn3/rzHhr5WQf0y/VQ5UuUj6WpmGJrrHCJzg3E2qXH
wh4zLKT9TXUknbzPxasNL5GLFut9tvUPb/k/SSISPGejfaDKtSQ7DhIi1jL+ScMP
PNwaXGx5o8HzCipFp3hha/3v1AixTfdzkia2vzgsDgBmgPSvNd3G3d8I9fU1j+/c
rOj+mL9SdpDhFTkoUj/oI6TkzmNLDSHNB1SB5I4KzR8rjG3GaYHUVhbWxbNfiYfL
JA5WN9lkpl0UeJEvhfwoMlA49lmQ5l2cQzMhy3EyRSo9vlJUjxXDFHJk4aU+O3+t
r8zDLnKywk9cpTZCgJHudqCtc9mNVhJFyYPAXerH/V9hv1bqcgoEBN3q76aIrFKB
LIzfxCTHi1aeGJGUnA0ohtBBF/eTZdaqDL1GfJgd/eggLUSkzzqrCmKGu/NrOM4G
VvFpc01a11JPiSyQC00iHqW1xiIe6FIu7EJfg44vZupl4hawIGcdu4gR3g0WROQM
9LylulEP86TpzowS8VEzHtlmNoQ/6WwytQJwHsOJMRnlssSnha/eJgwmr1shDNfR
l8hNHSzTYFaplqH33lBWzWh59E/B9t85YfncZ415gtUamROW0QDpmFY5nr/7eLwd
YozM3Bj5oNDArOzg8rA4uLaGZ5cWOjA9fVnHSXQeZWKxFqP7gI1LduHTSiR9MHZd
ru1ximOrwR20iKe7kFUsQk2QXXaihlzj3rn9Pvzw/ToCL4yLBGZb0yrPaF2tuT+L
eXlhBVVAB7LFXVFIWT3HhWNxN892f5yTmKyUFS3H45pVMsNGQWqsiywyAT3ngHvt
Oa/r/e+U3s06ALGPpV3midwhylJUnSZWGLBQ72452G/ynyTMMFgeH8itDr3ZqE2y
Uw4vo4mfnbYZzSsRK7wJYGT0VJ6moDwLOw1ukhZDgNmT2ihFyNlHVTdDil7cCNjn
dDgbICPXzs8HLtiUCQt50FxdhYikxX2EF6eQO4No/cmckNkUFZPbgt+NM27DXU3d
+8lQrh+YSBi6j0YWq3BRXZUZWZSPFfrL23mO0tBA3hYfCjgFnItfwy3ckRjVhTQ1
0ubZPjD4+rl/mZaePIcknnJjnOsI2krUtUhQpniO7ZlnV+DtVUktWj83fHMLqlvV
oemL5O0sA7zHcKVhv/PBNN8+rucXtTF6vk35yoMvmYt2G+wRICfnBgKzPsUkJjii
f9qrySTC5+N3u1n7gzGJTIJNMjTbsyOVj872tvcZt2BEz76eAOSaBRlGQ7N60J3K
mAJ97GMB4Dw45NPI4h0Rd9r6JOnXVcXoO8UJv5XoId23H1+tnt+XHxdnRI2GPsvl
F+IhxcFuXg1v7i0KoKWuXUYPy176Fa1u8hGct2Pm5R8ujp0mmfZ+F6u/FAVm+fJP
e5CelxUIehAPzyYt3+KFC3u0OojlB+zcnl0nE+7UvKfPDbj/trwGbVU31NntiOPZ
Rcp+ZUEHo+g2LC0ZNXQ0RVHW14JTGjgiSoWriydhrSiACONiVe6smGoi0PcZv6zb
paJ50TBCqtkoJlJuFtZdqT/hOIRrt6W+YidGxJyz8I4PCrsRCQXET2tXx82rf1vv
F4PuQB/4MXDmtPY1QbWRCtfzwv7a55Vaps1mNJEpKcMAnkz5f1bnzOn+42K/Syul
MnJB8CGs5WlJuxjEX7Wfxs8y2R6e1gKrh0zoLJcUH6FqLtH2Kdc/1EXoBb+3gWqC
TmPIEi9vgNrQBnzXbf32djtLaho6DN6F/ninS5oHw5KmLJ53yklsG4vDTSmWn9wI
ejk610VwPGjS70wI3rB2hnpk/XAc4Qg8QE1dUy/N5aFm1ElIhytjGDb8ShoF/gZk
C4cCYPT28mSscAlth4JRvik0R9RVrQ3njQFv3XlJJ6fqBSO0YCTcsgEPNiqcjAjT
DLd4yU7HXtQl34+FsyjwHEqg257ea9zURVFK8jwKCLhXA3dNK0wBQuWJ/jWjQOBx
pTFMvzD4c2AP1YAMTeWG3L3yxfX9hXfVOCH9GTjKB/pxCU4lRXxIZ4i3eaBhO0d2
nkBDOHZCTD2lNKFhWKbSy/zzb8fSz4Fir2iSI0Kw7gwx8LUt4HpQ/c+aouh3xQSm
da5SE37nuBtnQQ3KRpevvGbu7pEUoAzSbR9Fnqx/aDtNlW7P36KqVF8AdPmeZA6K
KWN+48C1SLIiFE+LdiTjjU96VzC2YLbrZxzlOenOr0Q9TfaHvJ9TnXp5GfH/M7t6
kTdo/uEd9rgc8l40i1soraArzysMoGdyaa8SHbkGFgmzM4kInjJlH6i5enSKr+JJ
Kefny5ARYAkKiXDZ9hqLXB+O3YUgnpcrDPPXJkB8yzwGMKHptymA6dLi5cV5ZH3v
W9LSfJo97JeoLEdzabUYSsWBam2KCh+ZNSXZdXMOACgNL/7VwY9REytwKAIrMpUa
TDWZR83CAoFDsV5uEE+DQqHTZ26S9gC95oqkamR9z/+xQIWL+ekucJcFh0I5toHj
Y7GJmB1ldZKrSOeZVNTw/AKPPRr7GGZPJnNOuqZ98qWxM5jRbzZj/xcl3V0/cGe+
PVK6eOcm2ubLK5uyCjHqvZHXsckPPSRnXYRWNoJ0VZzTJkiEGD0RH3AZLpOnSuR4
M7apoHcOhqXy5ARBHf9CNSMqcy9/G0zQIGc7/2eQu0ztgwLLYf2HeVMKjrUt5h9x
FldGPGfi4MhhezNibHcohem3rnxg0XV7IJGi1WaTj/STDBt8z3VHMpOONDX+bvXj
ZftvEo9IDLl0tS9l/nVNC77jHFJRv0FNFFbMvybqlYIDjMyBAryHWmqASxuxVx/7
budzZeTynpaZljfBVivBkgQc///FADFi73DricQf7+UgITmmAjxpFMtX8Zbn6XbN
DwxZER7YvEhFdzUUJd/gI97+UaGVjt/AxoYGHArl9yEbBwOq2Zt1636aD5byL9f6
Cd9dcNAsl/gLR3dsIEqsfGFY8CRhbeWsDM6WzsqTIP5BHfjAPYf8bR8hYBzFVPwM
DSZjiLqpu33+uAs/fHqNchxUZIeNmagvkPArqQGvmGs/tUPZyb6a3XKYVgFxyU2A
CwB0A2iGmXX6tCtpz6wK6n33/tFxuCSzexL3zn1/7pPTAV8Pm8jFjvb1w/5ifpNS
jLqB2sWLp6/oWlz4qupg+OAwiFDMh74AnGQzqpbmoOIPlYP4rhUhDd/MBqEnlyMJ
bcL3NltyUrEmYhhCdaQzTUfMqZ6ynqdSUx20jaMt0zjduDFrR1uy7IMaFRTyvQF+
mod3fDGlfqp8se+q3hP9oTMKf24ahb+62LXIc0+zrspgZdwrmemg4cikFEWUXYsS
+PVUtzSLaX0+WQHgxK57VuRF1P7C5A1XZLKdrYQggvTc6g2Yz6SYtYgGDSun5eVZ
jTyEPt3TQR3x4jTnk467l42rH4GJ+/0XlSnmUpdLLO5BJlBwx7+T8S+HmaBFZL6I
4zxT7LQSlWvYPrtgqry9DRDYBLQDvvgOWZ9AKKOB/M6CCdpllnlgL2D6uCygbnnD
EsZxnbz4YXDeFr0SYhVFx8YF06fKUxcnxcSSXsOb1IfWSj/49L48wcDXQ/hQ1Ezb
6VYwiKITvHAYt1eXGVenOVXefqodVxo6Lq2l+GWSpRlm+LDjP7evUITmfb6zMUOf
avyAA8eP1gFievDIHSKpMdulzJ24nn2utjh8nL+PkoTgxlyPtIRVnnI93asmuGou
FjfkEoyasWVewPO0uGT8mouxYlaS2/BfcVnXsg5C5Cs7hiUXNuISrMQSszla+jLm
uvutY7XgthWx7YPWu864XvxcsM21ikuLXDy+N6h8VZ4kU/8Y2r66WzWojMvztywV
HvAybiJvtMCstCs8SoQcfUyqgyX2COABbm3bquk43Bg3/y+7lAYBjjPZrOoIZWVy
7wVS4Hr1oX3d1/FTg8ewRI/GYEx52U/aMptEgaJtEceGSHkEe5ES4ZMF/buVSnBn
8Cu7z7snoqqjsuWNxVNnOGrFkCPcfni7X/j4p8qkB+UOcqRC4B1Tvj8sex+NmLLM
BnTPQT4RGJCEo85+ygYQdh+Cn4nH/2GmgkaXvSwpK7gIal/daPFxQQs58fxUeY9q
47TyKGhejxQcSv1LwKk01XGREFjjrXWoL/xGE6HUXE+twK6nt9O16J8zXZX65nhy
BvJF4lhb9WlH5UsNly8BFqz/gZ442P1DzYBgHKoYtLStBNLKZ6I6UGb1jBs805+q
8MPcticgi5zR+iZXhl4mAiKqcDyL+aCrMD4fTuHUEqTlK931q2ct980osaSJ926S
3uqhQg+rZcSceFJZBfosk0/Kt8yzTimVncoH1wWoHA+Sn438pJHVXGqTuAxppXF8
MVLdVgYQ8BgfhG94Lj4KkfAkW7BJ3ZCqzXE3k88jW5HjNE5Nz6HAU5mqFhODnqyF
7UdTyEk4IF6Gyxm4PdSMcy1T4AoAqtDvNFcLrnC3onAkwVrhaNXFzzdBjgKj7eHI
akuhSL2LF8U9sAHGJ8/7t4qkLgovzdAUmMkccN7Z7VLlwUhqEUEsn99aqzzuebP9
q2IqFRwcSo1XFJDVt7AcMHNBccZXv67Wwpmm94lcvsaCapygSn+sBxGsbP9r0Pm/
2fZcYZtp/C14sum8jrCyjFBmdTwGM/CrL0RcyZhEGPZ5iILFtqfgfhbiLIQ53S/O
shxSl/7XQoi4OQlDaiK365PTU7lzzQEf/A38A8ISrXeBXRbXkbdm5hVfUXgEJb4Z
6NuCRKObKmIjbEpQlZgygzu3YBi2EAPXnVPHKtkr7y97nu8Yxkgt3qDcGxXv+MgQ
9T8lj3J1Npq2sgpqRFRCPZfR5SpFHn8+bUYoC/CyuqrRzI8GptiA7CyMRDCDjwB7
QPk41ucEh0QM6wC44Gpopo6NcNF8CD6ekpKu2eaCFRKimyXMTKLhkCktQBMN73sv
WQcRLr1eca4iI/98e2WYgyA9vK+0A+bm9cpNpAMIyLVlBn6gV26vmsUVV6oKwyiV
jd5UV8CPzuV6OAlOaUyQBRSQySE2YOn+a8QJp4VOtMBL92iqGNuMX3ntmF8uWV0D
wVhMkJJkMo2zWwyOJOonCivrTC9EufPOhFZm6PteM2JgJ5ErdAroSt6C0zTEiLqR
MKngreKhSLxFmiUpufTeZ64nFj+A7woL82Q0558FpN022viMJUcUHWecUwxZXRD/
EVzoS2tOxoyLc9h2s+2TUkydbkdUk/kNI7CqHfko91vdXt4xy2aP5qu0qOlSJWX2
3os99qEUvFJp6mLIgFmmPg1GH8NzVGpINYuRxdrKiXqOPq+alX/AfM8MAIz9wxfy
5r5Pyefn5e+ylIGAHfy5mUwe24DqjfdKNCNsH/MOpak9bYIbXlfbM5wfdONRPeA3
JmV2fgLgaD/KxVGeM/vnQi73XwlDCdYvG4PocLNoUT1VvKrFpdB+LIPagJM7hbc0
wA2FEOb4vBukOfCVCk7X7aH19TxQA+2Z7wQEx3+ySqfFXtLfJx8K9OtHDIs+UNho
JCAkRnZeZxUAkjfo4Wn9dXZsJGtifswPMiE3DsouHjqWS1RiRoF38m03kGCMsBQN
+AJ3kuQ59yzFOjY7vhHgPXhqm5rSxktB7+9c5qy5+Lpps4cwZpG7cOllgiXzrIx7
dGdmbos80hsn+DqMmfVbnDFPJH2m8VVssltXfeGZ+rWixqGoQSQN1UbWlif/FbWc
Rg7YKqZn9PtMY7o32jN+W50Vpd7SsXiq4rAF9loLALiN7pcGLx03QTiO2C4lIaOR
CPhIL0FiLAtGUg9GOmeakwwVnkcW5kcDnYhWHGLmLpuTOG+wjXaKZ7kOc8BJgudx
mNxzt+JyzdEUEy/w1I7RXXfNC9CvbIJuW5X+MF1vaFyud7lQ++ywLox/gK8WYrLB
MpUw1c6Z8jrws2LmMHQJ32jO8SiagEVpsllPJg5LCUcSkC7e9/E6VToNgG0xeqEE
g8g+QkuiKk3Am9DQ8SeKq8zl2kL8WQKMC8xMyDDg3wBqkeklCUSEmiTFAKtD+SBM
dBerC1yC+5TKMqGQ6NZlx0dwIOhJtUDx1gwPuQ/w17u4Ze9ZW5ZXXv2uiu5j5pYa
ieNwd9lN4L3VtdmoIv9oYbxg+iU/dKEpuZCB7Iv9G5BO064769XdURtYygjhBiex
ghkQAfJhXqna9dPQbsCf2mmGF0Vgbho8JE2JUzLEeR2FnJMyQsC34FVbhHIVzkzS
NFxrXoiDMaeWmrYjxXuFWlxskj6ZaWdC8Q3zbKCbFLJh3QW+G1SnV57txgp2QJ+3
KwGcgH0YARGQmi9s7W9NRzh79MbHTLngmNoZwFA/GlbakFUTXH6N0lF1vKOfh8eI
3nh+tbhFo2bK4VjA+Dzfn6mMBOJS0/aYWUBBkn7+P7BoSwcsA5e9fyxUuK+wTx4f
NzZFCltF/V0/R06anMo9pLDJJgepOhixx4k0Om3mIeeQY6kTC1CIoIDiA6SyZJy/
PtuHTb+hD5Uj+crNOzsuTBqt64P1TxdSrnyN+rchYn/Hqt1mb6AO1lZcg1XNB1Sc
KpLX7oN89cyvJJLUVpVtqckIlqpDv9u+DZEiJt40x6xJRJkXsqi5+WiIlQK0ZE8x
+sKVmxAqdeETAICVmPYuokJGJ/cXO0LI/WD0O4CSymzpzzia2uD6ejTccROYFxYs
u7z5JVLarRKfcvtIp72AZUX8nbG5KBXaCGaHzksv7h/shmOjwLeO+S1n7UlNAbNo
6T7egUnojSEB7U9Q0gEbD5Iat3eE52+DUzgs/QEOOJG+8pqkvLmN9GtwssrWG8sY
6kOTNBRtPXLgrkGKErxXxKZCO7TRKHNYlqvB08enRqV8pcUZQrhGE8yWxaVrGQ9z
7FbhyN+tbdVd/unWD9jGONTUgeOLqQaD6Lp83JD45b34gDTo3haj7gMJ4VcexuMY
6kDg2G2P05zme2Xt/01x+E357DORS5wab783jg53rZNVO5HZps0zSCCHOmhNW2Tv
3ZyGsluPiq72/5qaefzA5mvpSXXWEvzMrXRW/aQMTLJZJ6EKqxUT6y105g5KBXLd
AML5tSz+nzN1tB/Xo4qJEo8v3v5eV/K1KytPoJsEmaeIK0U4kaY7MvIQ2hwhMRbw
/hAFKJOveOvTHw+JefzOCtzPDovS869s0FWPCZZFTVMHT1b1u49NmipCN1pafepo
TsjC4mUVeP0qpam0k/i/2omp8hnnE/cYIt62+ZFioLgr3yero3bGTNr3oiyOL4Vf
kGBGywFL4ri/mq9G0oBseq+BgRznStUAmQwzSQ1pcRYLu56quALm/ULNSqnaKL46
IJp4+IVBjCJp3723v3mI8h9BsJDmqx06rt1RPT6GndtL+ek0N5LXreykAWMy57cu
GGn5GSV3HxQD335TpUGhHMWWKcnRf2O7UAROpxxYExFVZ4fXNXgmFmonYHqTTyc3
sLg+KZAmbeoUOr3BWDoJVw46jTSzkhs9V6w2FT+ZSK899x62DdgHk82FK/UQkn85
hkPBdbcpY0BVpIF4kfecsOWd10i4Lq1QaWn68Y6p1Vhczl9sSh/RZv/5uBFVC3/9
/TqVVXfG6FFvG+b3ymT+VBcykWJJ06NHLhafkNRDaeyQDvwUxv6tyBk8CCgHl0vN
KkdQ2kXf8bs6driIkgCr5M0KRTsmiBIryuuNmfqWuEr+kYslN7q2TUah7TiOL5or
V0uoBAvJyfC6idXQxqPN4NYbQDQOd0+FiyOgtwWhqi8U1NBPF34PpnlsuXF47z09
TalWUmhU3B2gfYHOS+ZGjvpHU7ShGNS4EJo3jjxaEwKL8SkN3LGCby8lXLOLMaOq
u+eRb1yPqThtSvzi2v/IKhI5qEbMiyiAJxpcYQNrHA1XyAtfr48LwZIl5MA1WaEg
r8ci2NbWDyilvs1dFLI1fId984KaDmX4BmBSOEFQ5B69yG1uG/xjbPEdGTEAik+0
tJI+gcldTegJAf7p/+p2i6QOBJdDrWD2gxZg5qkZ4aDBFeyYGXh68zbQX+OOaUUg
aOcewiDrRcUF1UCqUngx9aj0o13kIOAXgVWR497aJIuRoDrk8LGaWn3ArLAKfLtz
RmZe623l8ayqee0MlEa+QMbpUPGEcYjsRuTlH/KRoP6BuZpw8YYesrhNe3pOEnD2
zGNj5ZF21Phs0BbZRl1z9SNwMSJO1VioGjAofrqEPpxxJ+hdlbr9AORN7WFZ9/zz
IB5lI2+1zD8WpfBZfFHgLuD42LDH2Ua/4Tx7XWXPbHqAf+94XHSB4kfQkcoVBnbD
794LHYAGGoySZHufoQjBzoAAA/6rRtxjbrPXKtFTrppMLJSlPJV2JAqgrEmdcL2Z
GEU22MCWNfAYL1efRSI35T528e8tkw/e1YXIhTJGr3RFQZdmVAihaI0nWdEZcPkk
e1mraC+m25RvHtLa//wxHc40aswrdOvMCK64v+xn5FU7cvy3Gh7BCyiqAE76cM1E
nnU1W7hVq/hfOA/XkazumLTdmoiJDd7QR6p/964j2pC8cDxJ4HuHWJ3pOTms13cn
Gmaq556PYZFKBgJWF2vVffUwsgHahLLthPpV+bCtR/w9a3sLOdxcoR1gS7XryvQ4
7GVgCcKBcn+afgyEDi3v+LriC38xVLotv7/O4vzNQAIlPJ0+8sM2XyallfOfhQPh
92HitvT/e63PjMVjNl69AWD8kcaG7WXwCpZEtCCn3M06o95rIIzZcahFAnaZFDlI
fxuEGZ10Kr+2GEvkPbMkCxBs0tzXTc5iCWI4PDqsTLK27fvFrlG4HTW5H11jtRx6
Ux96A+2Ht19OaJPGH1N6XC4IfHAnnwZsq5r6c91bd31bgUFreM11Qw9f6kPvwuzL
pRz1w3AjQe/H8RtoOs74WcDH60JOdraVR56J0T/QpFBlzqBKY2GJN7yqgCrHPUNJ
dpT9XFgXnVbai42OXTvHzIJlPHoz6/0FNfUwLjGT0yPYRUWBnsrmT3mqRpsPLf8Q
MxEqMtRrsMl6LdpF1xd1sm2geFsMsKTTdYgYxDPDti5LZjj6SUj+ISL0g8fP9+QF
zKwcLMH8G94AAzrnB/3ZfdB89bvz2KGR9Q5gGu2IYnQe48U79rgOpOT4X6kLr4G8
WM+Ibyujso65Eq+GXlXLgql/Sf9pEVHYca7l/+4io3xFQApG/wi0l4wA4KuD+WKz
jOEHB20deRvuo7MIRIMu5XCxE1V6IaODoaC2PtZbOPon77DJ9VtDu+RfQ5s/rBcX
Dgib9495l0rIofm+Yw/U5BrYc1aMJDA/2zO9+c5k120r1FyRE6X9VEc0IROV5+ih
yYCMFf2gY3AX6srZJSCH0kOqOVmzDvmEs/FZfTSnuAsgGI4ksQZ2QVMQzshihTSO
F6Zq2ezBcRbIN138MUSRghYqM4Co4ZpJxfbQrPciPuVgoDZNrIyebyPVPONYhGAZ
vOxYjue2/vKlBI54WEMATLhCSlqP3wRFoxgfr8QaiBBjDZf2iq61piIU+28ye6ew
9cQiXSYb0XUB+pFpOFtOij4d7lRTseAEoy+tFCuh5gJgw3ku7ZOvsWCkFa9oyWyr
GKcSyQgZT42jCOosKsqKcs3WWbVu+ZJioSjt/e5UIZoMfb0unHK9jzgih8deGHro
qHcEGsx2I97m1K7/FI2JWboZIb0Hu7xVrjSu6LixnJR/lnSH2izksnbiMlRvI7A6
YoVcr0RE05HAMeFqxLaC2LGc5BksQFrkP3m0ve2q1pGjMq37KvA1jeTat+GpCjrn
epFOUTv417rzyr65VMWNt6VNbun/jXv6GLZAxzMjJS0WtmW6pYmuhg/3s/j3iepJ
GQqX4YXown0jvBjhZy4u8db7LQCsBnNc0sdyvp5Tn9PqRYbDzi+PEJx8MXZ4kMjX
kv3xdqyb4is5OV/dQdNtLJJaAbJIhvy3oFLaCZ7MJMHHX5UuHnLZZw3QRgsUM0H8
oHFOoGQVlcQwI1Rx6GZkJps1n9Dcus9PFMFIrrgx3m6N5wkIzwPVbr9ShfFguFvg
h+k5EM6uAJV0g5ZGZK40/WzV1gj6W6zpZZNFBCJCY0Sl2iVlmJ02YA5GnDQFv0CE
7spRmO1Dqp6HvjUVmNMW6E5MA3ngLAV69sRv6cx6LAqf4vbWHLHhOtfCbzJZ10T5
aVfrmHwfNrJtAhxUUPd/2s0XHTstTx4e6I6ZS6tWL095FPVngy6vYCk9YoKMt3ox
LuHNfx+d+iHAMIv5UbYKUrGG5aUjxK3y1sKXhUaSpzvV4OYONHX+uN29LPHVBns1
XwptNXkMdEXCwcTp8E90RGbcB+C0pxk/UiYM/ENCCqnCBPJZou/veVCI0wuNM0ts
UrsgY9Ig1CPdJW0aMUqOPqcjqFT0cnofRP0XeKyydxandJnvSOxeeD8BfGT14UR5
PlvmheqdjQOmLP6DHVhzFSzSvaLzELrdfX2Zg8PRvuldmh30ujEOt6dh+vOo8DFx
aESYXT8fIPP7gluZ/N9ZHPgEWFWjRFxra6Msm2OoKYSomghQY02dJZFuO5fixEn+
ZfYSpcandZzS3r/guRcNWoxjpwyYFtq2UU2Xxlzb+XN3slZUl+TZ3mC0uMyu1gpr
TndshwZDMKUzVngIrjlEVl1ABvQNvZ8kX+p7LsO1UrSn1eKOc/7sko2xx69REcmC
CiovH6YSSmdFgjTk7BqxARiCXyQPjzyE0aMyfZkaRTcRnly3qP6RpphXuJBpLRH9
3zz1/jq0yksv1UCJgr8mQzijTPTbYuBgIMBpjtdzcbICm4R/nkDFKJYu8wLAlGO5
w00k0DAxwlceUBj/62m+nzYMDidojMFS6x+08p3M/i85rJZ2As/unO4PMkMfUQhA
8t++2HjQ/aAxRrGd8HKPgeDMpxS0PiSHxFDr+cdJGDbfXYuYVcwMn1fD+hdqddiX
CRTUSujPRGcZOZJkRVnAVzstYHe8miNebqHXQi2Uw1NMv4FC/z4HHj3gf5V/hfbW
1fvTlwXRPyVHEwylvq3fL80T/quYG5g5CizJr53exwllpMcrmYclISiSYKbHoMwV
jXueGEawHwohwuOp88j01V1DiZtE6DWp/dKYuE3MDavk+Kf0v+Kd+ksoPo/COBiT
GugLeqQ7pIQYPeHL11EjAw4JswG7GCUgPrUBot+mC6tuGLci1OJj22VXyc6Mo0sz
+J13Yk52KnFW7MQnUvunp4Fzr94MWYIUNygHtY4VFZsL1Oosl3JvJdSwP0MDN9bN
KJFLiskye+Sy5iwV6QKFGB8wezxEJKITMUHYK2wfwekvvloRoEWnFCGuvrENyR1G
NGAi+09WT25WQRYTrDgQAlNX4zJl25dYClm0srkE9hTH+ey2wP0t9+Yl2WV7juPy
oLlj7pK1WZgnbOBK2HJn9k6zrh0rHUtBWqhvHMTqMOFEHoWwo20g51VafZwIeBdq
foOMnjfbngjJCIco1vRGQ+3eR47IgeNyfmMrux8GqEbsu6XzzkdvQdvDndUXh0+5
9i+kDjwMoaWKt6Vhq9UCo/VTiBuhecauCz+Iwv21xP4IMSEtQk19mEL6F4Vjzf30
EEoyr+AGmgXlsx5S2mpoPwF1P4Ch/5Mlke6fzjUfRmly6KhfjZNZRnrj7uuQGb8d
BBiANfA5SssxkQzPXByGaUkSKaZ8c9IjCHeb2wkAtUQHi1WfA+n0MotBgkHiWACW
Jz4whIRi8tFD0jboK8HHt9kobHcjCOagvqh+atJSrFqS00qwuz/wRhykAwzwkdg0
24kqgKr0qPKLHB31/MVXx4QblefMgPyMAgujxmWYEfHXNQqCovGNUagJpJXkC+64
Vm9JTF1IYqHVNxxBYr+nnGtSbbFU+G9JJ+wg9+HYwviXIRCQ+T8hEE/Ml4OKnDqI
a+7PFzgyuNphcks0A8QvSmgZ/T3m5NrulRRCYfsxBPWeIcBiRnYH0bvrxtAgSaBj
/MfG/hUJPLo+HF84RvsxzrT7AtFpakOwZYWflnGyAiXgEC3TkLdPESNkPO98WkPD
hPvxAJ6GuCR3PXVBFgkj7rPaOlfztrbEpYmtVsro4Mr0j/SxwJwXJobecOWCcpao
AXQP5+2TwBVtNRAr7MsDrkQ+reiBtgAVgXNBk7ODNQd4qUIcE0ZYHp6gykrKssL7
tk6pFdpTGTF13q4ygwZxSg3QDrZY2nn/AqwQjcp0QbtlY9whKiBnZGrc6pU+LQeh
ph7mFjql8nDWQ4hEWxk9istGFvAt8U8LZLjErYQiD7vv3pibHz83u20/HmhPpFO5
jO6hNycA67ujc5UgD7SYjm7xZriAIzFpmfSwZITXlgenIRUojlvAfkEzqtH1dJkS
nyBW/W4nhLNeKTxMQqHdQiAgw9w8s0Fe/B1wVDwbyiS9jj1oZH+hN/hMLSAryXHh
3XoQP0dZWje0xY13wk1CIJi4VPkknXLbr4ID3l8kcYYbKej55d+0F6tXRKFiP+fh
4iCRP4RnhGxjrkhWB87ieUeHqP8+LpH4H91KQl64dgwJi0hSYPYriVEJQdIw4QTq
KF9fsLIqBuO6RtKYyX3oRc5tXhSR0F8KDZ9BEpkjSiftU9uyUxE4PS/EM0aMM1iB
ZOSTlgEJIis/080gFq7+vqwZpOMk0usLKMbbYv/HrPzk+tUe23p7wIV5FHZPhDcU
83YfNskGzsLKnFkoV1hCHKtybhhRXEW1wdoJRfPOQf73HScga4LQIHF4fho+Plxl
3DI7QQpCTnJmqq79wdNPooZppXLjt1y7Z3ahMYCSde1I11D6TqlJgnzNn7+YCMgy
bhjKj22/NO440HEM47Kd7krM1rnzry7IKG4KqzeoGZQRxIlJTg27pyBDi0BRNRRj
ntM+gFQRb5aW0K2oJxivZu1rZHv7KlViPdRa+i4qUohCpkIMcoqjjnABOOHZoyuh
VqiXfdLE3UFrwmLJGy6Vh8vlBxpJUcHhq/h9XVEaghL+xMAr/OgD8YvV8NlJ1WK8
Rn6z8LBXsISf7pRqOghj2aOzQehVxdDwjBAtozCWnPYEluX6pM/lbSp/e6qBMkGg
WLOyc/Wn5ieqzAI4IqYzIgq+94oBe9dvpvrr+WS/HJaQaibadAv9vabDIWTciKGY
P8re2THwUAZdDzlLExkJqNsoVVSsX++cxZ29sZnXu28aI4WXi2pdkWhZaeoMHry4
78eCA+CxmaC7aEFVfNMkUgE2Hi0DekB7Q85bBk5ldECjJ9VZBcWx72JSy1/xPbDV
/tdI1wx/WtFjv0TFtxhxgDHEYCilSB8HcKNkTFx28izQH2yIIm75QGdWF899RYwq
yGfMAwHRcGeaXf0ftBUo4SMb9Ta254mTsXlktLZQydY4YbffnNU0Kl2agxeXSyVN
QB0w64DxBLzLGC/wpr9TblYY2QBds403Cq3upM9DRr4h40nHv2eEiBqddyUbTw+a
hEjrPnERhjM5FKiEOm0HTfsW1sc8mrB+wW1Lfy1SLVVcEIl7c/fMmHR2J3DJHfLG
u8Zq9TcMfo55z8pDSjrsYomlCQg8k2F9nQnTgjTc84lTtMbka0MNhbB4FvdDMEkT
UBaoV+2/obtM6mdvxeLO9YSxqW9IVGrVVhvK91S4pmX86a8zYsRuw/MSZxdrM/pC
S5I1RayS45P2f0852o1//v5/bVW0aatiypA6Xq9zf445VuGpaYw/OpEVvB9WzF0T
kG51OJuv3u0XezOa25Wyug/uDLCfcdMqLyOPc1B2wP6CyTjbEaONFyCOUFyvgUiH
ofp52O70oFMey1gPlTBjoSV8O7yDSznDVIt3NYgBFm0KU0JXtAc91PmGiOSlIu1i
VhZyCRILP8A4AJXhLlYA07IramF2iJOItUkZe9t2zKiKYVsBgQZ1ZrSgaQFWfK6y
aPR6MomHxGzZDlVoh79Cbb/J31DHzU4ATDM7Nah9Fnq9TmuDPD3cQvXsbUFH6qqJ
5Du6UXpzQ1rniS3kdWuxzbYZOPz4U2QDNC/39+JmuMnVq6aEbk7Qm7YHq8PInMQa
UOze+V1XWYwxZkBqP/u2yu08JYv1W038Sq7YUc2O2JsRApFcK/5zczvulHy7QIGp
vxHclt5v4DrKzABi4Ow8m+4R879CcuSMF6eie0Dz1/+icDkZJ+LkTFttQsiKDw6+
9fQcdkHcauEXD9LsMUhQ0E3PfByxMhVInvwFBRYVopPlWLpta+N7tKAmTYyiloeK
BGIeEJZ0x2k3/wp76DAAH2T7O4hLgAuaZxmeCir6uZDi0tzBOvK4TG1kLkSmUSUf
moslxqvRTCWm78p3U+2WSrWwEHyUa5PQJ65t75/LRlAQGr1X9zcM7zuPdSOj61WZ
N4ZmtW/gFXXLpuJL+7AJUpALB0yiFl7hfU4eTPvdYWPQpyd4gSbF5cb88xFbI/qS
yw9yIMRuH/VJGx+F6/KJeYN2GZk+B58bSSFka3+Mr2sIQtb8+EjqftC+RcE87e1V
Ek1OBNnTRv8wbRbTKA3FBx2TUq39mk1mF9ouE/J3/a0UPlBqna+w4fvsA48+3aQr
8B1BLqnbPL2TJCWkYkOGDfgjF04CJ/cgKIUUHLkW2xTOrAZfvRb+Sd13JASK5MRs
dQVF9xNqM7ZKGQXr64Am9384DtO2He1o4ZxvIiJxsuorEyqlgXSoVB2co9oqQN9n
Zm8gSlIq1nONJ1SYqq72ZKgQ+HinniBjpcTTOvl7/hpvLlv5j8bMuN3yTt7eeoRn
wtA5iWClkUPwz59gzpUeqe/RimYd7nRTgoRInWm24BBEQfnUtZ4IUsi+BkjVKuqZ
ighWU4+qxlACkjLOooDBBt0yiHOL4aylnhiJolEfPr/I71O/ysWmyhQpqRzLpxtO
G1SDoGoBI1Hs+w06c4A3XwleO7myxDF/xIT2qbc6eUutRwVTw21roAA9tYUnC4HE
xQVxZcuCJa27MmR5QWx5fif9yxzegN4+2jRhj0mh9ZrwF0A/b9s2We7ESJ4WKX44
+uFMttug9pz3Y65xa/TQEK+XrBBrCdfjWYyHkKuE5qHGKwR9Rwr7lRYjXKFL+scF
iCVH9OJuc8mpPLAqW9qRxE3UawIpMYH5HYWtqv80mfOXf42mgeDuHQpuXWJLPFce
k4Fpdn6fhdIrpSTNW2uGat1TqWEqbYcSlhd7+Gr1mT8dv8L91cWcj3FZqWUdnjpf
11zv71P4V+DOMXBWNjLktInZKkwRoUM8p2O+qbsb+f72V8SuiibuTeexaHz9rpYT
ImZbHznFbuecNwA97W+En48c74tL0mR9tNwzXYInbknDcQg2yNnnE8VeVtl3kVLF
gJsGrroBlqmArX4oJtkrS9Hr0aOLK/wugd04BegKucFLAhRfXSiJA+qgqnq+0mux
SM4P0zdsp1jNA2VG5c0lyGRQSBqnKwxOj0JzfHD/iC3K3g7xeTsBHg/cvqm72qBh
PGunx6VvMdOH/jOM8OSHBVMRWhg5fCnt8H3mvYdzKLebNApDNtIrPe3Yhoi220HK
KTMei0UXCl9bGIcobvwIsv0c9pHs5J7d4/dagBnL0XdqBCYSeanJZ0YkSI5nwWqN
4iOScEG+BTbPpKIKiJOcfAiXBkd59MxaDejWaMSH5x/ZURBAjQ8+UlfRlky+hd1Y
ZgrjmeTVorIxe2fxbqSsDym/JVL02kmxGzwbtTEo/RPlKQlRZ7c4oPdbCbe5ZAPV
mF5u1XU1DNAsCWb5LxvPyxgeZVr3vP1cM+Qk0F2hdH23bdRIJl23z2ibny6QsRS4
sl8qQyGSyL2R4gGmGAyRV8FyNQMvvnTl/ZdLc+mr5wAtpizVGKmScYxJxYdRCOcj
J1HDv5D5u/cVYDFB35LW62+9QO0zCQkvJC+o79Y/GLUlR9U1HdJajgaBN7LQhi8p
NyG9Fp5wGSUgFKditwR/YcOKffrdOofX087uoQ+0Ofk4tOXLeGvRKbsnHd0kCBIO
FhGCgsWyVpp7i+Ocf7p+pWru9K0rhqYd70WebqRSxSFS3dRJJ8pHseaxajl5ur1u
CRrWRwvqpXpyhEAI7CMGN/KNTlIUakhYyBXWiPf6gg+6sCk7K28OGB9z2UYk/bzx
0gbhQRLtBiyB11x+6JzdqJClZrfz6cXOX7CLGANe7w8AqI93CWhYaMQc9THOqlxC
dd+KPf0st1keo1SlJFVxr/Lq7jlkxgobr/wG9ONGce5sUnqRRINaZqgOO/oOQE8Q
R/87G89G7QzCBcNfLSlWG/tMOh6swMi6kiXkCAMhwMcalRXrFD7TjMZ1ixJREI8L
0aH0j5ytyLRhADPcWT6zsVOW6w78+iYsmZIymPZYpr2LqgILORMWMkAehP/QOMfp
5x2PdJIX2J4dNjLnPhPKZzFRlX8rDe37I1jLqIl8euaiVTGQWlzHHBP/H4ATEt0t
kyyiKt7mN8FtBeIsc4mhCFJqDdp0rQ/rtOmGZYUcYCPxMNuAjUwVPU+NvyFuTVeF
iZJobjnhlW8DghZq1Abi95XlK5uU+5Y+2eYboaP2Q2Qgn6FAIWvb3PGlZsjzaM6J
7Lr+6C26VrK+8bzMQdKAQ1lbz2P6uy8+7bu1ecb+5Hnop6Os1mes2m4MxTp9oo2c
zdWwVUqcQNV6rBkW0QvEdqvK2w2jCOHzILTfIlltn9BY2uaolkrZ3XYH1wDU0n5U
XukwkUWyGKVyDzryQx220KleXxAlh5m5eL6Uthxcf93Y3s4EnxZgR/2RlKD9TWTo
ByAW9Ocj9KK/vDvujWnE3qb7IWKdK5sI57nQmIp12jVKYVjQQeM04a80SGw8Vklq
QhxvrFQ/zCcAsTzZbTobasEl+WowsLASA+4nQfyCBkApVsea/LRUKdmuTf306SgP
QZSooV1RChiDpQZsNW+7iccURTHZZ8MGSiiXQlgteuTIgTed10rbmCCdJbXA8msj
dw4N7l1JgRBG+H79OJbJ+Dj4Wz9lsAjl14ucYN+VTgXQr0hMJGQm4XC7U8h6bQ+Y
8b2l/b4+bOx4nMxxj/Qk3qFkNh57N3OeNOlx4QaxwMd0r8+CQ3jVmLZhA+yLTPKP
6JRJa/UknEpqX2On8L4Q3yYq3IR1bLfAQRA+GTZNB9otAac8aZ745D0Yan/xUqru
Z/5to8a0mUy5DexPp5UhMHCASS1eNKioOUN7mPPeyuemr5QUo+p/H1aTr+nmmAXx
vfm3+CYG3MLSHMYpF9snPbJMA3U46ZCulqEjA04WM/ZwQourtb/WfgkGkt268/Q/
tIrWHaqE8fuSphuicm/ZDiLPipHApsoz2mx94rEwnceW8e4DwkyiJaUg3V1X0MvP
eF8CA/y5Unu2PTYl9ZuUDrdWpDbkNoL/SRQhcvf1Q0Wqx3ZDoxMNr3VgdLTnjYoN
SlMkv2sp4OgqEN2AJREUWPxaLwT30NJMwfz1T5bPVkLs+MYV3UqsaHj70bYHvv+H
3EP6ein2/VAzYSdgm657+acwx/PpiQYweK0CzjOg/jEbgDJblqlJkMVTWvfvvDt1
cETYqTC52a66ImzFby+w/HJnum5bT3beKcviWsGWmpK9NIXGP+DmXm/C8G67ygmF
hE2SCVYI1UFbEPAO5M+eEBRAu9BD+OFlIXi9GAGCnZbJa9OYQCZeP/NaOHBb/pga
cnOGuqq8xm7VOqETzbeujeIMiR1O9q0KEbIcmoMx41/Zn7g5rcfV9HIYjGWK04rs
FIL663cQTFW2/HJkbYRyjuijedVKIvvGQmGk+pcYcHJFTMtHjjsMZYJDrtvrx/RQ
FAdMgxNYLX6DcQCW43lS1FizYNsVF0NxNVjXXTusDBSQ3s5KFPlcoCmgoh7LXZVt
o+ii37ZtgDGcet85RTHHaZLje5tu7joTVbSslBZz2byHJ9AvQfc/v45FuSjsNtD7
9B1JvKRRqWAmldmAzXl1OEKgdjQj8J/2p88/B0e2qVsXKgGv5yYPo5+Vj0DJdLCg
e3cUgiVSzVszwi1kF6Cs9anNsejaSHN2VtPLN16ME1xGVr/1BRsRIy/l38GidB4/
jZUqeVnIMXdfsVf6zTxpCg64k4VTNqJ35RXYrzxhhgpSdw1aQkTnN3PuAeOGBaWN
lkfCuv6bvVKKFkQZCi7+mxC7eZ21t3Z0LHccvsYQ6ReuKt/qozXGAjcuAD4FN1KV
QwWloWK8S3MTAHXSblWdxrz5J9+8xW3yxqKp8OEGSgzuDaNEzOn1sFKXhMVcUN6G
MsMw4hTI5zrb0RiHUskjYyPl66Bv98+65N834QIEVHB+xzrVcamLaYT26C5ZrQm0
+s6rGMtwbCo8FqdFogxZFq7Z5phFmFfXWxlzwWRb7zh8F2OMc+gEKnhFB8FTNnIR
YzHosSaFqFHKeYZkR/JTK4SerPKrTlWgcC+pEQNGV07SJ+6BFvRmtNpDgDZFnBOT
DyzU8Ehh+Dvj+XtsJL3N+3xgN92WYW3rZNr45YvRIqodGNJYpKoRiac6cFJIlB88
R1RMUumKpP18pcuFZ3wb3TRyH9yryeop+Uyqk9xXqg1dL+mDhjhQzOBd5qZXfaZI
3zzcGkWqHxqt5rOdYAl+FXHUJmHV6BceaS9osH8/FVfS+qj3dxeAIIPVMpr5JW9Z
0Y8fA7pIgNrLUjRY9UiUEfYUeedBseFUkwYIs2EL1Uzs4suvthFVBeBlbYCCUqer
UK8mBy5sIMGmF6pMfftKGg7A0tSJ5rP1zKMVaQ+eH1fyiT8jbdqHqOiAxCzqW5iE
zi/YHGUjrCIYwJdTxrufUjpgMbQb4brHURM2jZr5y+ZlMy5amIPDpiUkAwQUbLI5
zTsRFZ2DC487R/FFAMJFXsrRVVG/jrv9DL5V4KypXuqDnqFrgx7+ZVwKYYxFx4No
y5nnKI5gHESGnLPqyGeekJoRg52CbprMEIls2Q/eXZFuO7ccBd2uPgxVG2tHXF6I
AnxK+vMAa3YbQlKcfm8nI0dj+Tewn7BjrWaAm16+w+iccFlCKvGll7QatVokj/Vh
KyVze3Ez3BP/EjuYlzBAyeAE2ixgQNV5OObiWt7Va2EaanjrKlkitEY8Sh+1dX7d
daQTa5JlIjBYsWe5C7HGr/O1HdELX3fd9wsoV8G+goqVGDEmsZzJdXvbe7UCZKWv
wt9pE29YjwG+0sF6kfJUUme+QOU5D6ew9ckGbwDEC7acAhfhYOtzxHqaEUfIdmA5
mWfwKwM8iaqTLVZ/aHzPl50a9uiVIQu4VKRtWuxkFmRaSEZHBGAObRBnafeAncXi
demZjmGgFw5rnaWxB5O8+BKPQldIMJ/mvm3cdSgTas0fP9EmzHtjPBPRDrMgdd7O
TYy132CYagaB37ZJyYHeo80UGYKIksKXdiABkL1pqnyyGEP7RZhU9DoySXkPdWJ4
HFtlwKDwf+/Qax0JALUkVyME+/m6MFzUhIkt44mGy35V41IK+ltCMcphHkxTgbJv
8MD5+x2BLolrgdrkKJ2+xP7VKb7Ur/PqLN9E5x1koiCKHCCU6nloFn5DtzhgRRHU
dk2CZidp3kZ2cu4K1yLn00nkeA50bQPwj8EhY53VSWSrU1TzdslS+dL5ameS6Nuq
WGI6tgPVc0lHjluJbKeeTK7jbKVCm8RIOEKcqqS+rlvt5rScRgbsXoifE7Fur98m
VCk3F+KALibj9VMAiN4hk2qgtxPMQMXi9Y22TZi4p5Dr6KsUWXxSbRPixdHQZSuK
kALBOg8lIW7TuPOH7ZKr0so/T6i4aQ+7/1kyJE8s6EECrWn995EqbkrEHmGKt3Qn
d1Cb6DekrsPskD7QoxI0mGNt/XhrM1JQ+knAIxcCuR7fX7k4QXEfmKdD5GeafRsp
QyfXwAs+kHMAsNbs5NWOJwhDyKRyihkmUkKzJnNMmjsWWAiSdOcbgkyr/OXZp02i
z3HhokdaNeIpqqv0TRsTJJThiT1C1ObiBEzevzwA+QxPyYWf7ms/L5TdH7N8vdJ3
rVmhWyveg14BbLyJ+VeEAHtWZr+HjCMvPyHcdnkjjp7NUXrF/Za5k8YfxvIQafNY
V+/02jKtQnAdytoQZa002xnlLLhlMfN/s+mAyU1YuC9vhQSZN2FaTMB4jnTOaco8
KsKHWCvI9XWBSXyWwkHtpYljF3iXA3Ogq+rmE5phvvkx/DQ6Q6riEEZlMkl8+vXL
8Bcd1UTsoVBdccxo3KekAXIui/j6L/nQ6Kw35AYQ98fAlaXe/oFCT1AO/nzNHxAY
aoYLO/ZYWabwtKhVREDmKl1jNeFnCDoMwDmyPcLFUADFGEdZBQwg9nzYXNJ5LlH3
qr3rBk/7k6tXaZeqN4qkrrsszBAHITPjMwsUcYfmeUd9xkR8NEGvI1nV4r/1qVLP
3VJqNCr6VZGa0JxIyYGR8JLZ64kdAyUB0pNzV+slf4eY5LkRM50+jl9gILy3XBZ/
B9j9V6yFMikM9t5u6gyKwQvvnGXrmUzh9qpyTL/fnErht+BWneBwSrxICbyMOb3c
63ZfS/v7X4pb1aVj54ooGo9sXtu2MX4m4qp0BUTYi+qyEBM3gxo2maufl34DQuNw
wiN7cedDyHnKO0LtYtyTUrmFi4mEkyJiMNVQ3AkNz5/l/nnwTZL5R71Al32YwOa7
I+Ldk9+9ESEZYjjGd66Wb0Ft9Zkrw+EwtGYAGT45lLYesGXx7tDDZE/6ESnT8saP
jNRIDRo+uJMRqZmjowF1qi0LW2eyRbwrdPEbgw4czBG1jHS4Nq6AKvJ3VqIDNwlL
16EtTn8aP5c1Oq8ypB1NOv+glF6BHBMolFlR7opCqdYrAHixzq6dDMMWOj5mm/Cx
mxMdmS4ABMEh1jxrgX9f2uy3U8EcfZNettKwIQFINOgTdtSnEOP0UeREbPeMlZAs
7SwvA6/ny207IweJ6vTzIyJ90/6qWfOJGRwbvNfrpV4nzFYGCzFSV7nU4lBcs3sG
hmUj5pzTD+/xeU/8+wUKG4GHK15w6bB2Q78ahJMZod4xzIsx2nrlSd3IJUsqeet1
7LryXGWfnZmLe+zuCl4wWN4SrAPLyZaBSBGSErWl3a0gwVZnxTun8jdIYKp3FvPy
D6DZwCBlaEajcTMho9Xmi+WUTwpDlkuhFe8LGeJNN1sgqin40AziRjoKcP/NJoY4
1GM+fOoRbMnEDMUVasca8cKvUrG58qlCX9PJiVpTrbfj8FtXDmpGNhl/IkgtUNEI
tqmzvKBU3kGSV22aViJ6z5LJ1u4RIlDLJQpsi4X2UgzVtNWpoiZF91xmgEKqCUmN
zEoYG7x6V7KZKVIPlaysvhxgNhnFjE4j80+2g5Y3TvEcT045Icz7LHS/hxtJAYc+
HVynA+k8BCD7kX2ZOzxpRe8U5NT+1nglMvO4BSMcBxxhldIG0JVXvZHVd/KXkTQH
i7VosCJ3hZTvJr9kPev1amRHYsg4z7TObwGiA6nk1VbVR9YUi1Zkhc6rYndIJnTo
3mGWBhoawKcDdB/IFtplxMlThIQO9kLb69afayOHC/d3Jx+71QunfeGmC8WAtzHI
7BoxC8UFOP6yuFrkb40nhtY6K9BXrQt9kzP+PHk5JtRnC5UciE/NRrUSyCTPphxP
an0Uer63rzzGZP86wJ77mvYiJ5cVYpjjfThb8WXXmKlCBKvsanLPQEeZyYcGKljM
yZdg36GI9LOIJmWmdyUf2CdfRe/CRBR8LUyoZRum027kHcamXJtqEZRENgOBBjCv
smYkknt4OdC/ysfTV7u4ZCZAlZVy+i8rC1LNgHsCa+0yhaNsWyZmhF8x5x2SEfXC
TFRjoy8eMB/wTDsRgI2nKj7hy5+ELYwLqFXW1jth9LP7WqcuhX1nO/aVG2qvd9+z
4TiFAnC15gXcEg1tLxgxCk3+eYn2fOK1frZaAHnw1+z8eyjMlFBcisAZte5N3Wd0
wXIu2nUGvx8H5gsvXIaVrHXhljt8F1A+hoRvY1oJLJkECH1Gxecp/YIziKJfXpAd
jG5ry1FgeZ1/y9cE1dfS/BDGODD+7/rthBviiPIZgWwilos2JsbfgDPcuPNRLLjr
tQPt7TMOy5EZnO9MXk27TDAqJ+aczB9cm2RIN0CELBZyw+f4sd2nSEhg/ptEwnjt
4/Hdn0qo68gn492Ni6LO0dsLdkJMqu/l+ceySYoqLAqPQ6kvT+VJyZkOCnHofaxC
o8MScZAAN5vFUra103rUgn/cvKcCqPG+XML+7DIffMBQArmCzTWr314kgiWAdUW4
0uAxtDWWE7TEqn+Is0P5K1oJtLMxn2QsVQzcgX8t0ppbQEm9sXlvLI1seFaekciu
+bO7JYNllMEo91RPAaggaY23Uk2tnaFGx/9KXZqOdqagQXJ3riiQv3w776L1I9Cc
568jSKKsW4jQYC9AEDVzI/Yy/uQHZklnshMRQmvgluUXi0CybI4Ww9Ef8WZPzO0t
nexmdqIWNYd/MbHwKwWjxj8mo8DYnOCDOsZzZQCqxgCCnIOMFyoAqUotX+Acb4bY
R2teAeFC5rdbQJhlU8kjOGuGR7xgb8zPs6N5wRlxrn3jU/ItVYEJzQhQgjFrbpI1
0WCnGlkekJNSvUBraVKSfr/ahWTRR+st+WPjyXD9oqwlvrtI+DW2nF7w7LLIWneV
zC5i/fbd6wsK71YvjLN82d7qaYdlGyaEuN7HZj0m+k02nA4BTNDHgfYEKnfOFzL/
dHPFDvBLz9mbpFGxae9koL6VhhJgCbSiTAbav7im8Xk7xvr1qx7ElZFLFNU+gv9M
nrJymgwDGnwoWeCA8wuGL3vtLH9l1Qzf5dm4r2vuLBX3V7QprWOrwxL1NYZLltN7
ElIoOX+ZHv4oT2nAithL81kvMmF1S9Bcv+JgVOmaIOor7VBVJY882mM64OI1FQYk
6kmnlM8k3jOUtcPxvQwR+l4ETqVx49NUrxd583KeShVirEC1awiuELSJkDPrWCJK
ivwYqMgIf68faLMjKeXO5jLDwjH+04m6JA759WgKBdY0mSCPOAsns3526TPto9bG
W0StKvne1PkLHVIH8PCvGQFRGxpIuiRdLScFGMGqM+8OBe5Su56SRWiVxzrAc4Wy
DhH4MJ4/yf2+JZRDA7U3vv2XzoYk5UIg6DjQmjoZVxcBoJPm+1l9Byy40Ms/tiTD
ud1NUzRRruN3nTLcMYC3GND3F6Mgd0QmmJOnrjrPVD+TibEfzdocrvGegs3rm8Cv
iHeuiqGDZalyT5JoUQ3bNButiU8jkDClbXOKeUUPLC6CDVCWFTQFqS2zegluBohs
Ir10vpbC9hh5f3DdQW8ZwlhBBfBXfODJGXF9vnqw/ZTS9s/v4AXb+sCJbgxsmLl8
rPUNK/Q6AXvidAZCvIk6Dtq32e3DBvrwg/OK0fMr/6LnlCuRvDgPDqpGELGIHAS2
o2t5RcSHbSGLB1MDG5Aai5RJ+DBu7nkwUeMXc4aBwpc7HLEVxaQRLPxBZqWt4vIv
alNzozlSJFLhfntyk7xmN8iUKK+wb+Y494zv7IlS9ohYivHG5Qo8Fm6Tj0OeUMve
OuLNg+SGUgJNrHStis+iZUF2VtQQ43pRpeNjmdcRO+8NVjZU67CQpAFLWAdGk6c1
Z63knWEyoswQd76O0FWtkBcGQvXXCCndHhirtqzAbDHpFA0F5cB/FjYj6+XvVRUG
lWUoqxDUF2xCxhtQtJ8zPDe22fxMGdk1VxMnjk5+dhCAys0+6+gKPJV6XPqukx9K
1XTO0p+GtdXl03/C6p9eUdyLYTkFbr8QJs3nXhHBgJJDi+3gdj6s8++WjyT9sUsq
FMENIkXYAEsR60TB6iUkt+qS4FcLFmTwOc4jwBNDktTi5ZK76C4He0jCxhOAaJNu
PUVxI+adrBlnSL+a5uwMfry5wiwNWdhmiUkMXGGtNhFg1OmNO9ACs0X4YmbqVWwz
sqBZnu8cTr74wf+C9xx0lPz5PifPFEvjUGEmZpu0QbTgb/4bJbOgOV/911hL5H+Z
NcaiFO15890xtBpeegS/fg0ivhfvKm82E541B5U51IgEJQstqZ1H8+Y/UThKhIXo
lxNbeH145AtX+fufMcrwTlg3STA9yFIpYc5EY+GksHF+g4EsVBgNTjL85LIW6sk6
cJXN9Ma8q7zqnNhdXFuwnPMRf9FISWuUEqdmFwzgFDnoDVYsuozlUN6bvUA0fD2Z
3NPVQU3/ONFa3pESGQAyb/v6bo8bNQ8aDR/7sczAqUVzQGswJPc6bgtGIZKse3hv
gXUQ9c8EOih0xbIZpXuiHHNR6LHw+chKhD0i3iGSchEy7F4yAMGrdxtd1ZBdb5Wg
731oI7vjM9kODxF0onAI+pOP418soQViGd8wvn4Kvyk3m3msA6/1b++LJ+uik5pS
PsKbjlkUB7ogRY5w6lNa6/kbCm0JDSeWCP0CDZHoYvhyhykcLHawTd2PLmXg2Lvv
uoNsY3GM7dZpNbt1wry4xBIPsgqQPHdtp45mRYWsPnVvzKnG9waTBDxU9XjN2Pnx
sL8BgbmOYXjsAtfHb4/9A33UIuKskCfi8bEZDDzZqLub0jitgLMoOzB31bsZWm+7
mEljx0LginGgC4ylbAY3gC2PHmnclGAbiuQ/DmOVYQIHvHjzMSzz8TLJd6rduY0g
UGFzZ2UhfOis26L55bg5EjtsqckmsozMYJf2Gw1yzFTekFO34UQPmYWe76ajsyZl
dIj2Ua2c7fcT7gNVv2qAl7DSpjCkknS/qwsTJjkBzGITuWgQCK5qOPpgIFwiZNGo
y2Zt916hWY1MHCzcleVWBtjz1W0XWRuU+Ad15a9GrAximR5UOAt8k78FExkgzrA+
IZ4UeUdANtTtIVt5iz5uFo9VU3F7/TkMX0It1USed0jsKvrGJLCcOWxuFuI9EqrN
adlSq9xZuLNKUt7v7KLfNoVbGJ1666zEgPaGwzn4xjFHHxHYJZE09DvYWJgjAdLL
deyRoje5IhFmhoRNHxC87++j2y1CSEH5jn9kFYcdTrDk8LIuD1R5jYFeC/gEv49R
sAP/jLBzNhGO+o5vcqZe89ipsAPkMMzbmQnA3y0+EVR2py9JX9xp1DajGD8lhHaD
iCryZDGVF0mpedECe4Nk1gGqff4zPcq2gNN4l5djWL541kYwe4e4D5og7Vwoo8rL
2jCijDllfqELi8kZzOfqkvsA9oQAW0H14RuvpkqbtrqTEN0gXvn4bI2DzuER0Pjw
8Ztlon9IrPEQ4GYy1yriaVt/vmwm1nYGD1Nhq6T9U/4sVSIikSn/koDzJZVOY1Jz
lf/VL/8BtPUFZ8Vpe6su2EbqzYVWetbg3C4v8mWB3xdstSxRYzJJiT3gIsVajz2d
W7eiGcLuIc/XyX2KEsVru7o8rvI3iGf+zMtphgPOVC9hjprmHVw5or/2XwvmUf/N
vRHpElpvaYg4G7kcDD2PtaaSJKxgAFYS9dsm19Z2mDh3KBIdU3GuT39HlXXxW6NL
QOZmHYFyJY5/mcnrf8hi/l4XHtjRPc2Em7ld6UozzZwx8jxPhpw0kGW0NGwxlrz4
pWhTb8BOsK5YSIj+T6BRJ2FwJ1bGXpRqaoohkKlJxwbVnkAEt2ayD9s19AVxzJRW
Klz+FvYYptJZQrouX6dWkBxAEBMDukoATVevR9MhESf08Vm0tHc0gBACvxs2LkMU
49gf7l19Y/4Dm9qxnPwQ/+4NpU83o3BLkVk9CXbeQxiEK/bNCEIkGL7uWyjRgR/0
9A1CyZ3S8hJc5aKAddsP/XwnkoKkHZWD47pAj0z0AQPFhsiRxEyiIBZcNnCdY6/N
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
AqlJcBN35zru1sigFEaEMkGDmuzpoSNiY/N735r+ppZS26haqY1ggncXhDrmSnoN
AXXicfqsG7wqfdYsarzIs6HLqNj+vobbBe5PkWguGkzEmO8+WieNa52sjkw/1aNe
ZAihhYxdvbxz9apE/DlGPMkKxF3J87mUXwkuvOK9XzU8Q8mo2ClhIfcODSgnfKSh
fCCT7RjWvO/0sFghxfT2uOOqkvEwoPGqhIL9lH3r+wS7j97op8PNt/zoXHlKGDBF
iZbwa5ZQIUZyl35ybFl6SUrqJha6XirOaWjT7pmcM8+IfONn2xyrVEEqMyDnbq2L
8qkwa93TmRDbQqIlmYXY0A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10032 )
`pragma protect data_block
r1B05345IX4tasTM9jd+/bYbCmYfcfnG2jScJPF3vK7UnBKEawydfWDf1nESP2se
Ncz2odNFxozYNOiDTXGpVAX+h0Xn1dgFW4Os1dY4al0YYmg3nI0HUNmGL/GjZ8N5
fOsc0XkWaoO7WdwDIuefpXhQM9dYfFzIQ+e+4v9hncAKR9HLKUIwp05fyuDIBUqM
sMnpJYInHuCampmUsPWr3OK95PI2pOyGikSItE+T6qHvMmbz7H+jsxnb9uQh8mn/
d/QzP68TVcWu5dBunnS3nzD8kXBk+gGv9ni2JkZvzw0OnD04B+pbUyXKmkYXzZ6F
6M4+rpxdmKvoifKUHgKf1KzSJ5fCZ+jvJeyp+uumKhkojMC3NRKXSNVSkZPBxPch
/usDmvGPXXhqqgGxjSOtWGYH1Jskbpiv/qV1p9D+qYZtXmYLJt7L2tp8dRmS1ASE
dY4KfMnIQ/zejNEEhDMOh4YXL9+Y/Bks3U+QAA4WicTzVuivux5FKB93coD8FP7l
GEPK7tz5Wzk+D1fkZTFZ+XTC+uTJ3RzF4p5HEZKbE3AgcsRQJQMseZlmxWzf4gL/
+PFe2FoMDMsvnQXYrTUOWfi2hk99dHqikasNL78BpvgN/8UIqpU+exDRQSseIbhZ
z+NKYDln3pdnMb0qBeNnff88DXo3oFi3MF0SS7N6KCPKsc4dopT31Wta40CkPT+v
Icc/0E2WQBsNbPo89l82b/yR9RGWsDEwJ0Q8wG7VdKuwKv3UlNW03xbKMo/0MrJm
tvk1vILKYvz+MbsFZKr60doPcRM3AyBmc+ctpwASUbjWz5+hO1PBRO9FpGa/2kxq
0gU1cnOrlOu0kDJZ+u8Pc/IuNttjIbiCjcRIZnp2HZvZuItcSjNkP8VCz3ICjev4
FqThm9cncJ+B2S8BMk09i8Pox3uouaAtmiOqROFKysej1l2efYdj04LaZNAjmRP9
PVI7h1sNtoby/HOqustjqrcF0QyvEvcIVYA0E5qg+r8OOuHrxcFJIWd9gZH3DE4H
KcSlwblo2WntN4IovLmp9Q8QHoT1j4QKyXeWnDi7/TtFf/cgb+5ODUXUaZ6sykka
mv1QypfClewuDKVJCfJ6576ezJE3dVvXfjDKhXzMtbPI7kyxMDK82K1VbNS+a/HL
QOrM1FVsxo9eXOypzRYcjleaGdgvZL0PPMOYBQvll/aHCEjaARlIA/Zdnrd0NDGl
qedYtUQ5s5Q5ZHwcayTAhbl3l2+BLB/E8hLSpdJv2/mUndidFMlx5u0eNUSgzjJV
4GZxBdo9msuhUhvQ9SuXcbWq2kR1idIdj3JCw9Q3vmFVMiryTRgHD66UYZ/JMHaI
bjZgg1Mzu5lt2IaB8yg2QzRZUFblbm7DTElkzUXtkbpjEdTQZNBZG590GC9pQ/ZV
v801tJvW9vgGNwYW0HqTJljSz5Oio9i7/xDTKWPA1XJ/nvoAC0RT9W9phPsEWcT7
2lWS5PrOQ02H80m5tYUc1/sTzoKOU5QZ+edG436MxZDrH6D0nENFemfbYmAXm01X
+/qaPQXPPLFpxKlnA7m9gmtS93miXr32cq/6iJsSTf9hXk3XrfgfwOK9cILX1WmU
E1q502WpAvzS0PwjYRn6ajiI7UqqDe/PMV4Z2MhBCHTph+SZWuH7nSjTLH9NbzQ2
LFeKmsI3l6pHjD5Ubz1ooJnvjipyDq0vOCv/03vmnc+S42v2yrxsLEDqwojuhJld
+hOxTRfTIUERQgBo9QkMedwCkiihRBhbLgJRbAT50A4b0EC0dZsg0bEhlK57szIB
aCIL7LWw9+nTnEvQ8nNSRwk53SyTE112wV6Mr2eT+oGLSS3XmDIcoMNoL32QdGlE
U1Ib9OSwB/Qrv7733CdAePZve0KgcMbkhIvhM1EM/GdfR+XfDX8ZXQw71cXMm34K
p+ZfHwkupha4/XDxl8mDJP2H1ONeTsc1krE5ATDvRR+Fu3u6Vlmw6J1lnyO6zrYW
DbpGqpgQuAcBAdmHJLpo4iCuL2HwAgxP2ZZ3IV+6hdcDkNaPMvlMMfrYC0/qFy15
OMTbXALukBmb8lN5DxBTNnjL5OzN0eDCcK9mqFIx9M3TvOi0f27hYrgKBTa2OpKq
4axdRXGxqbr+sckPbd7h6bzhjf2iEAChHJ5rAbRHN0nJreI2sIjRNeFqgr1wITLv
SLUtnQLUA3QZzEN+8kp7E8Wx72hM8d+hh/uR9FfXFTVJavqRtYcQHQwRA9DCtOQP
RwA5i6LJy1Ob9h526Jv4NsAx7KCYTKfATW55ga0Kv/FjaYa0+0dadk7orIxVny+Q
AhsIzvAinoPTjw5Ac0RIgPPvWyso6kDi2aHiAXX+qcPc1W6kIpwHuyrQXkk1sr9K
mPv0OYaQUTxol/6+EV8a5Dwf9q4SczgtsKP0pBWh5MyNh9rJh0BY2k9oCBP+Oa2n
pQwgRaphF1KVTmP3vXZ7aEa48wMrHrPDJqCTtbajDHDp5Y5fCZ9VRoozcM22NU/1
IT9fQj7GTswmf7JzSyr3oQth8KMi96UyAeYFUeHYVro3Q4M3FbCot/bNhYIhFmq7
j4q9gOK4Erzsvm8wwvPVi9Vy/7FWpHTdZJJrg1lOpxwISLkwkHBfEoE0wmxICAei
QGkglULOU5IFzlTfcIKO7AAgSdNxbtplY95+IZswoDSyIMBVvjGjuJFq4HpxJFOi
S5o0H//MLx2qcInnYuS/mXmWkH5mXTdEHCe9+tnUWbMV5V8qQXsYBOksxpN4a0aR
1fEcP/N3Wg3P2+x31Un5rEhxUbVv2s29P6LXUozOVruWOEk9CkNu+eUtZcRQOTgl
uh5uuZF1WDjaJc0Pqve5zlvewZQWHDccqfZDF+LbGSwiFI/zQUmAHoiXAj6Z8y0R
cK5ZdzuNaNm9wsa4cZJGgDSonZwOqA2f3iL9irNavZkiRiWu4XAAIiiZd0jDJlI/
DZnL0DU997VKdO5Pwms56SFklGOFMarApsJ5OQozxUAaC+vWyFvMs0xigWoUAWjC
luhbAegu3Tw0S7GJYb1KpNK3zrdpDnYxTuwXoTz1N3hqssjPxtF3bSjIN8qdu56f
9ZZl+M15ZDzOLeLaoF/oge9MR4wqqaFJp5ohLFknl+QyvcSaBfLr48drb5B4B9IH
FnxxbUIkjR0NoUWu4TkebGYRXm1ZwgwyiwZDpWEvpNL5b4UZ21Ig+P+R2hE0K1/0
aKPh9LXoe30khkoM+E4/uBv69IH6yX+e3SVK3fcj/hCFmzgZIDIgsVJVUTzqo6yi
I5zIwBu1K5BBF3wAjYsNUQW+u/sUFIIdr37aG9fvclcMTiZLLxEUxd3TOri9jexp
sO52/YLdpx2n5uQRZN/K9He+vdhnV3uN574+gnsJ6PCMNPolgOsAwy/aiuoP25wd
cK2OM3ocq0XXYbpQVPhAomrbB97p1OXWY1jSrhgv2nwcEv0/57YxtrnlgxnWdxaL
ZklnYAYmk3sfSv40433V9qrhS2rYO8tfmNyrAWRd1Id0IVxbHvy6dwpI7sZ9aUg6
C/N7rs0jApjgOKGiFCoG85N3YfnjbMXrZn4j5tlgM1RbdPbk4smqF+6wwAm2FW8j
EhGION88kfGV/NJb+hl95iWZacDEWValNbzK0H+ja/SVBkyW/hYP7K+hGvkpx+fV
wDq5OjAHSi1rphTxE11v6Pryc3/YsLF/qNqrgCdpc1T+WSXasXbUBn0h5otf3Uzv
/TEUz1LGscfHZIdn3tPb6/WLzg/1mMLmfzeixRZMezelu4+qlouBvXq8NoLKY9/N
OXo3EQS4cH/af44usPIg1yrH4sY61LYDQi8xoPAe9vjaaRgcw4g5iIMY2Xy3QTIV
/FbEXTDdJ5F3JEcnKp0FbwCpWahYuFaHrRSDgH54bDKcn0RiYzzLNDWW6yrZ0adt
F4X9JTAvLCchQ6GV+7pFNGQeXiVmaYd2kVYnAuaeeII9AVEo2nc2zHuK1q/qDneC
UXgVC/d74/9sMA7wPkQmIHEQQaSorLqB7yUwzq+E5DJqlfNwe5hiJz9PE6gVkDjJ
t2gFsvINLcn9DEAzzX112pMo4aJ1HLUVwHFR99JuPHGTlVXzwZ4RTd9y3OlfeH6i
dgQuuMmdfdfJ1Figrb/fjstBn1OPzAoPLo586DiDrk8+4PVuNhPJD/Cvn9nT8/Lz
0OPPaOzbr/LhxOELl+avzeDcoj41QabahmusG9uZWTCLTWaj1YJ2TJK02iJBW2Kb
sMchB+6YxsWQi+7oCylpKXfC3TGw2OapZ9ugoDq15tWiTYFk3ZiSxKkO22KSbUSj
BppYI5Np5PCBBZWy/SWtz0IwXdnIMCUorjWLm+kScUEzpOSQVPw1haQ1JWD19I5n
r5g6jh1o04k0i0nskfJ+XEduXVfE9LdSVeAcGkMjhXOPhAlLLQkhrlG0minwKFal
lTAJO4hH3UOHcVULHPpZJft0Kg2voGtww5DDkhKZjTNs4SYMrXMz5dSzjwwVneyF
kTstPv4D2qyO0PUEnAICs8jGTxUNE+pniNGYMgmUb48ZBKmqIzSQQqnUEuEmAiXF
ChAS+7IIcWirWJC4w1tMey4qkElb7S7CeyEtdS9koHMBmmMr33S2VJrq5KZ4AQsA
vlxOe9eHpd5Eb0T7OSXc69l/zH78N4DmrcSMZDfyUnKAqZu2WBjoeZGK0jxNlc7O
4t/ZmRFvlQlBpq9UVo42s4UCkQknxuykZu6W+gKqCKhWJvVQVwd/S4nviuZ29TJ3
buOvWP/uboc3ceV77yqpEm99/uXCna/MwfjtgPESiJywbi0dl8sPmDGtezMDXoKr
6Fy5T+ZwpY3L6rG8OICbMWIzeNJAx5UvgJc0RK30aPnvh739nUQe1fZS0FdsIUEV
WyA95AX6UmLLJfvzu/QJkYHwijk/y/Mvezsks8TgiSncMZg9KljT31KKmLXA7d8J
t9/mEDc4Hx3Vzfnw353dmPWDblsUMo9dpeYk1RrLBSJco7G7sEpg54dxfynCSC/q
X47Fx2DIGgSwK9BfhhMy8sFVGCqWpa+Frl7ZjyWvN6cfX1bamoQxa6BkkcLd+l1p
OiPG8Wh1Q0KDiUQfFnz/3qIgB2rAh8CH9Ahps9XxUv2TEhygDFb7XdRKhuoAKkzi
Pgd4YKRNSRvbeIU3eWknzaxWAQBeIvuDXt5a+J7ANBRHr0ErnQO20Mt3sMo/DuTZ
MW1yk8wxSsxV/KmQeYpyk3UnN+7mNLkz01iofYOJ6iKWNn5W647Vv798LR1bzwcQ
9Pgko94L7FulVQ+vK1D48RDZt3eTiJNGcoSiDbOWR0uCj8Uh61IRXp2HrhIlpccz
TkNz8tta7Bp7iil7f5CtHKeaawW06iymPi+04VW3QihhOMtCVKjeB8HN3c0jdWXc
AwnEtBIlf67kzauVGntERDvze0oMS2HyCtNi++6tiTM6dytrSPQJT9HPQ6xmA4eO
40rD0OitnO96mmST8uCR3u6MzTwdGNHCJGu2eXsygviVi5o1uKhh3NaUmGyD/hCu
M9tKZ/Y/XTCXPn3maBl0NjQ1Zb+zup1YpgbR9w6KHlzFrvNKTSnfHuFsAJGH5BXg
AXp/LTQ4nq4QlzdrT38vA05TIZ+inqbLl5+gB6FWNUEoSvNxxSXcrYM3Pi4EZUSv
mS8tV6sc/0fiJD0y1o81eyw2jkFN9pm+Vgm3zDVNnBmqXKnxm78O/FJdbUCmHAWI
M0YVg6X9HVwgYob3WNv1vM6TWJmOEmCkRdPLLogKn7pkq7erzrxJoVjDqM3gc9Ex
XBkIa9eqwjEZKWBkNH09OhvuhlzUPiFDSUsg9GcgdeCBE11t+K4mEN6/bClOFGHn
wtzwflvxueLrFht82WUQvApkWwQerDb2cnuajek4Q8Ewfpquw4dv2Cn4E0X/aeZA
tqNEmuAkrPFTEBHSafGsucLla00iYuqEy3tdpM8LGWSfATB/Sm21rTlZbhCM92Oo
9QYu+j+BiNq8Bx2x3wo7Vl6PvFGhYGc7iDsxTKz9zcaYO4XPNRXKVgI0bsjO1Wp0
7gGO5O4EvXjtw/MTfYh+bz8y/F9fOV416E5QorcB2UeJ6H7IboscRl9oazTabjkn
oiGSIGyjG4TN1a7046N38KKgvzgf74CdZAiVppLBBtBi35293uD3E7SsDgiWxDZj
AobIlLy6jGYhR8r8frP1Z2fV/A57bAqG7x9olFjTYeghS6n8zaJaWicE81ty6BZJ
LU9p6bcPLB/IEVwsLhw3Of4KhdG1OFDDXtvgWYpy+/5fQeRvYzFdDyOWhlm/vNlk
jdP1QP3vJ+uhHVCf0d6G8DGmE5RtV5BRHouVvvH6U8+4J+EhTlISwVSzJMMSZwNB
jquG++e3lvqT8gJRSBFcrVb1qAkktWgIScFu53ZlLnY0+Um5Te3JeQ9F3YR0euZx
E/LoOWv9j8o+7EwAbVtohvD6dALDs/5kwqNLLAFnYFkx/hXD8TvtvHwfV7cMyEt5
GZJkBS/Vf+pZVDj0WnD/dRfG0MuesxCKIe7k4wIq6z6uk+lYFqYkEl+IRZ+3OsGO
ad77TkUJAAtdOha9yl/5oV04UPfRIUJutZot+t66444CNw6dyWorFG4Dwkf9ZoXb
VRNtQ0NvPJBRO+snvlQOrBBeDtAdukZo9zusbyrXNiZzJOqFLfKL6fQuhsmhJpEf
vCad5+dApos1AVrLnH7hkc8CbLn2CU8mLWSvOrQlbzXNxx06ys4oiQhhRbEXrk9Q
xWtWBkrCUaflG+FSEdr6XDFGScBSZBVRqkrLj26oAn6AiJD7TqZOMwy0vW8LGvsD
7t03b0ztTrvASIVbYnLXzSiQbWnTcPLTOM2b3/BklJAhsOJLGyXrAbsNaF201iu/
EfUxVUubiU9pR3Kb9IZKfb1Qs89cbkJ1ShhrJZ3PBszqmHDtSXt3buN0KkQBD0kX
mQg2b5k5Jg35BEP9wU8enO7IaWPfF3H2ko37nUe0mWGRfyg35xCO169YO0kOpzov
UxewVEcGE8h87CajaSDJhNVJi0bUalDnJqBjYbVWnDMGjdQRJOf87/s3yQWg+Ega
B7poYhdO2/yLroPUMJw7PHwO3EAUB6nvd30Qds2B2Z3vDacERJ/z0jatLEL0SP0p
3W8D9M5nbw/yFA4dOaB+54LKFtIRTSyu+JeNbEwC0oRfSYFJl9hcfk4u/RT5T5xt
6LxASZwpevo30lkz2LMZimfVIrj/Hfm2f+8Zy9uPiWCtSAivnRnQ1lSechihPNyJ
UyPFRaXw1gXHxtANrNbWMjvl3FHocdLlVMEXJfR3gdYdWxfXsTMM3fP0+t3ynufX
Qo35BTDOL7S0T93j+Lqer4Y/QNa5OrGgOcaBcGL7pqEHoB4DFYHZRTbtDiC+cmY+
/yW0Taa5cRWS8EiDwCHPp5QC84c/Rv7bNL3pCGUGg8Fb+9NxXvrwYiurs1Dl3Dfz
1CyWTasWTRTmClyK6ZqZEZ3gJbx7F/Yxiz73AiI7YdeJ4aQbUbrrhybZ9rGN09P6
8TPY9nkEiRN9aWicraqxMJXaf1igv1GGZ1pTEM1BTzu7R8BKtq3VDV8AfyJHUejB
VmQpmDMorY8nScrt++VZ0EbAKN61WAkHzYjxuTKFIGOLmEMQiMIP/naRfx4Y6MgL
oB2QIVfbiKH0+mmRY+t5DQ58vNl5ujx695foAHzLCQ+lUfjWbMgS5n9bnCAvjLBk
FRBIUq3vZUb6dJvVVgF4ezH19AeFU3fpVrNB6ky0XtsEjruXSfU6/SiuJI6RNyjG
C4hcXz6yW8x+Z1qP/QuBvPYU69i5pI1oVnHcI0avMgdsecCuhEQRmd91F6+fWGvT
7UzWtkttwGIpwWVUeIf5iAMC5kzAoJ2Xm2YHVAjXXzjsNoZZf3UjPbmTyY896WUH
ObmBA08VS2PC6x9gUKWO13p7y3HlyyCORrnv1/KJxzFu2bJIWIrQvg6o4mSBciwP
sfu7SSW5QNqH4VUIgcRn0GSPQJkaF6/Koejj7vO2z7BLbWIxlY08LQ7+kwX3UXU8
dWsH5fOtulVp/armvP5dRfUDZZdgoqso7g7tAXDVfUYIL2+rOWOATUjYCWgqaD/Z
/GSypCNyIHhLbPN3vW0OYoxHXkXGQJdfXFwYXDW/2pOnkE9SNm/js75dxkU7Kcbu
XZHdYlxVI+4LBKmiBpDxxFixb3hhjsgYCTvcB1QAUXbBgf9bQqnkpN+l0j3CkihK
luaf+UrCE4t0XLekYgIPjSsy0cc5ZOg6qw/QBitkg6dvETTthXxBnXlYjM2rCoB/
salt/hpS6U22WppprwoyNYZW//+7CJkGrp59+lJIIUqEYPqRuFNvGcUz+GuKMgIw
G1X13uUsWcyphF0X1FfCOTg+S53JRazUPfF6jpLdfoz6rbLrRYOUw5YdWWNs/6/i
6qEWIXmnlUwhEnm6zqJJdG3/zg+99+kMvCZqNkuWBZqJXjLBCGFbhaD4cwnv1FRF
O33xcBHz/u8fJcT+V/dcdKH5RglwO33yuZDc0IKb7tFNccnh7TYLXfm+jvHgK29E
yp37TnnO1IQKzIvCwFC8GoGEV+eoEMUldDw9A4f/vZuXfnxEEH+2YfQ1P657mwln
vvXIv+hk52WjaVYVYxXriSQuZ7Gg9jN0jkfLy8lpTFmD5l5AvYk5W+fAKFA8TznH
4XsG7SDZA2R0q4ynMY6+zjqc+UjrwKOS0up7i6Ul1xrmDa64FeScvNqUMJCHDBzR
oWoq+eF61U+NK+1fndiTWJL7Tnkl5qs9qRqdQMrpRlB1vqJXu4qdPqTyhxNP/ssK
PIGY/ikkbNEle+h6VjDYtDkwfmIbCmKzMYKV1XfTEHv00ucA4EGWXCv/6Yo0ZZll
zMKXNrl+UjddN9g/R8goASXWnK0kKlNv3TNDNbydOQjqTJx4B+gsFS+IzZ2mapLl
9RuJc8dnCEqTuPLE5dSkGmnu41enHp+ldNRT52lsAr9H5bOJolHBjKyw770XuJS4
21eGLrtjvAzDleHvnqpI2iB/zUmSJ5ZQDp+SDNJL5TK71bZ24nSXe0dhcH0RwMDH
NNWqjvljl53Z7Fg/V5nHfSRSs0VlnIMLu/HSxqtDsU/sZXuM4MFI0B5DgXehWhyU
OeL4fYlQumCv8D4uROH9qtaN1k+mlhjbHMN1mqiNOz7nHQQZdSryyOdbmqElHCOJ
VA9aS1ZeyFdCVLQTYBuIjH01SMgENbh5EoJdlvEnXVfyWqeMp05uyUzWG4EYi0x5
ZnkHYfI5OpQooFX5oOtiQrHp0ftyC7s7v48a1dnKXa66cz4dEIybs3SsxpKlMiNd
i6x1MNqX0LQRcbqNLpGsB4k2NVdxQgVqvn0kvzsr3e1XZk+0Z6/kphzEdJs3W+Yw
ILGz5HKSTbM+MpyXpW6xVl/E91X0wwHtioSPhC62WHwZuMpfouwKZ6joNvWiNPGN
gyqHHUrLk4KYPRiMKh5JbTqLEfvUTDXdMu9wTawQYQGJFZ3ckTcLNpacAkf87dPn
9h/qa4u65oR2UX9T/5Cd9Y6YEU9AEfGsvcafikxFawpWV8//IA1rsr5EmNcxq229
bJZPjbDQJg6LO3wsgzfut5zd4ik2Tb3cLD/9zYJexy3YvWnjhANaYhQaKQJbiHM0
9yYXR+BDAKHy8SlRcRoBngJkCjH0UhXpMgkfEjQdrYnY0eiDO53IgvTfWQ2gAigG
8HaNCn/o+pL8On5g7PsKl2Cb6vsVz4byvBppRu9+1TdBhNtwFX/SOrTmD7fLn5fy
auvAOkv0WhcE34VELBN0gue/J36vF5MKNmZcLJM8D2qhkXwMbpSLQPKDyIQvm9bu
nfOx88RTnejLg3gFo2SxleEfuuD8A27fylCXNidQz9PfN/TC46zxruktkB0GENvd
+ZcZwB1hHDNY++uQNKs3byFWVpZC0rRUmHo/D2hIWh8pEMZck4lxhY9hTTqbnXlh
3dgFSwIBm4/7cF6Mv51pnx0KQiIC4TeE3SvEncu+mOoBaw/8LGzgOJvJqJSOx4x2
UJ8qLFWrSSdcOy5krabtaWBY8j3ydi/gFAWTYo/xRNq19BYSHTJOl7pDovQE9Kmj
JjB6ScZeBhZw2VDOUIAoWUJWAi+sKE8v/Uqj3pwkZcty9JEKnpJPUCfkeNAT2Mcp
C6YYJFAKsJ47AEwcAz1tL6oSL6emOkA1OovMztqbWj5cQUNWzShavtCbDNh25SD5
Zk4Ns2TACkkSdWC871gm2KOJnNWHvNARXrSLm6eNRYwgafjcYqYzlRQJa2t3Q4hX
Hwd6xuRYQygwdpAmTIltMLVfgm8F4bBHXSkQlsAJe3FFExuo+9eoogru9SHwlr+g
sKRkV8wr0xVhp3DczXMmMj4oTgdb/RVDZcMb88ak+u0fcNSvH+ckgcy5lnW8GwKR
UvbsE/lK3rEe1yoC33Vrv+7Yv7qSOqQZE//wWhWcDkLdUVLbrUBVAvk2fIce0pXa
S4dJxbu+iXE8bK/sPnern8TUnApuykz12kCzl+eqE/RLgSzFqYG8CRERpd7LSZXV
yQRZTkrVWNUGm/L+OpPpIRTQTsvUIuyQaQTEjVIJdwMWPaVu5Zt3t9WMFsTFtKGT
1imBydIsHT8lkAKbD4GjQkyHts4Zsx3X5mRzbof2USkA9IKodhw+iKVVhoJjwdO5
iKqLxHaYBBx/6MS2jVAGayEVtw7yRpSMfAjsoAwBXfJQgcHRvJn4T/VVwV3NAOgc
As6uCir1iPLKr4nWkxybREhGwRApoKlbMbDZFROi+jVfl4SFYxyeW8NYkTg5Gy8E
4T3MbiDhGNOmoJgaRF35ySL78jl/5Z0lSZ5eh4e6rNw5UKsnSYvuBRB2HZNH6vSr
el+4O4dadM8ZkO+Y9f3zfn0vhBo+IqwIWR9eS7C47Wr8/Tles4YMtgJKxOPJKcdZ
/+4hHHd/zAdl8S6T0la4+wk6ep4Ctft3s9gEHrPxYK1kBpYV5EMh4GVzchly+15w
1CayJDerRaTPL9tpwaE5zrNvTfv9nCSBNS1f/rBz27ySBTdUpWlxQs0XWd79buPS
wDMM/dVSvCWgJEr3Ea5W8OPWRH0ZZnTubsDG+qQXoLQOwXVYoDyuQpcopQ2s5iqJ
KibOXzjhQTMZZYFxZ/HvPvVHZDfonrAVTDyBNWxa5EjU0TBJEG4612GCtJw3dkik
E8uUzCHM4gU1FBqQwxCaW76UFYbTw9ARWj7FxcNIPUWc6HJyxN3Q/qdq5CFTi8Mh
aLwOA8fLBp1TqKUXFAbEe8k8Bd39/0mfp001vQRm0E0wMdQAaHV9ju0v7IYiAa5b
rEpVNaJbC16y4gqDRizD9DQuumffg+aa8oXtHjHKAuTkCCbLwNEzOOkKUb+D8s6Y
nE3RShoByZBblqs5v8I1wgHTz/1CKuBHDNxmYMMBIvhGU94K0nY5eKeOOtV2ayIE
iBBy8mUwdpo+jGBxJhpV62SuZcP8HRBtm+l04wvCAEC4S1BigmLfRBLIMa33SDwH
Ku4452FjxW5TJOp5LU7sK9EppXykPVouza6xKmh3oJ8/EUSDw6hB0FSnl31a9Ml6
tHSPYgQemB4uVm9VLyX4rZxR51yEZnOZ0g9vrmIStKv0/gqmW60vK/bNExF8Z2Kc
c7PR3y+cj9g/mbPh0IeLZEWDODMgLwymLfi2BrQV5A2RyzW256vYfMVI79cTzbs1
fCl6lj9h5MU3Gwf3har2sQ3kcRi4NHu8irS3/cMBWIYyaWIuviklRU2roOQ8luP2
7vz4bGULrJMIznvgnlKbM2EkXRiwf+KkS5Bar6+HP32T34zPSEz2CR3PJuN/xldZ
ZJRmGETqX1FeguSgG3wBhfS3V4Yg2KcFPPyVfIVtQqclU8clxCoYogFBET5xXwsq
IAr0Pn2IHH5P2pQay4aC+JtPK+3G/XC1qGBtsCCL2o+AZCVnETFyE68oAfFQ0wjD
gvgag630/HKB3RxUdOATzrVB49pNWaMvZBLW3B3pXmU2lhAc8hdYKMeVj4v1tB5P
3VizP5jVR8DPXef17foLTxTvWZWZj7qj113KsHE5ijJO9vDPGRBzDzNL3mT+Lfbw
4QGEhjNaiT68a4oKpX8aG96Yc2c+eLEAZYMxDl1yg5sKauFSPpV04Qmu5Of5cpwV
EFvEIwwLCzURQ+Gleg9oAb9urTziA/bisVk/gpBHmhsyTva7/ChB2rfDeNlgUix+
DmOctpUQikLRVfmVLp5HfGFw62QVoKsxgto6h5+pf7ICKNgxJfmepEgercFNbYzD
B5QKiQ1mVUJGpnypp7kK9aIX9G/6DSaEgCvOSAcpabZGD8kNViDvgIIdaNNaROvB
5ANNJ0qZb9XkQBhpwH1pEXEzunwO10eEblxLXPpaKv0KKTch4zxvFUSoX7O/ZXRQ
1ZxLHSa9rrJr3jRGKfylBuprwG/38rcH8SAXFZmoKnjMfMhOB7V3JUPVe5sfGimm
MdwN08QEK+brAhl7S1vBPyYOquXaNeU4vk7U9lVDdvDyvMG4fzJuUlpV6Ddv0K4+
XNf5uHgiTAqbWmbNsxnqgH5WHEQfBYjKcAZtnk6uYaYm7b4+0L9BFLcGGZW9T9z2
uGEWZviUx0WHTq56DoD/ujmh7ss0o9u7q5jNjWI58YTAv775kwE66TlvGM/Cuhfp
LBgGPjSxkkD4XHOrDe08XGd7bT4jgUKnNcBY2cqR5PkOftwRLDzzKkEPrAyJy8QW
wJ5ziecgtIgmxFvypbdfPe6x3LbfHrIBb0VwlKLG+pf9eLk+aVCgBL4sLKIjMZ4V
qoxuNdPIwNvnCb2aThIJVpQYClyBHsztiNY/GuFEB5FUgVxYYafQ+WYPFxZG7ff5
04bdPCyaqddp/tegnd3hzE3K1RhNlDtT+7dXMeP3faqs7pTz3w4SsEMEeLGF62J2
YXRAZRzhdmNJtQ1A70zk7IksNOqAABrcCGa/qhWjBhr377IxP3NQfIdGR221+qZM
v0Y/eOwAKAp21Ft/fg/Ff+q1zy7t7betya5GIkTW/UvGjsRcp7kBmni3Iigz1n+i
Bjhumoa1WzLleLc7448K7uGqg1IBoDcsU9pjsZafY1zSIVXn7wy9Gi5/H5ihobl8
I+dx+VWSlm3tJt2/zbigV+HCiNUjYUrVV+PUgo+bDgBW9M/RdFYp9r3W1VAxo02e
YBdXQjdYQ7pXrR3YtwLTFjAnMAWtYASldbvSzMB38nfBLaBR3royv+CqWCgZSjaj
pIgGJ1pCFoW0afT+JRohGvAajvzc7qHiLglemm//x9/K9yUJPLCuHb8Ig322litS
TLtggyMN8huX3p8H77xPiV8UeS5sGx2UkpUlq1xi/hHpflA1hDF4nGA4onS5SD+a
RnybMj6ptgA2PC9+EzPNIFVzlQ6z8g3cJ2LyqHKqIBMKGlai6BUTHpeyOMTbyYTZ
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dl0dNBKxWlQXLpx5HopuhFkTWbrDxx96eMdFpsJGEJFBOEh0zf6zSvHMLgS6woAe
YaUK+APCfyj1zjkDKrP1OkX84xj+dZ69+KMAwkeH6nU6UdXDOXwgwVFtnSiNGGwK
I5Z0msZQ7uyQTYsXp70xj5guaAVCE32Z7QpLfmuedust0Q4+RcSaJpBFDkAkNwuq
UdCJxJsiLWAXzQhPRk6JAkMp3rLu+ZkJ0uTD48ypVvDElMyD3QRZZPhRfR2FwWLA
FaEcLvLbaL2waK47WjMglf0mqbmdVxVYEO+xXDMwgq9k3JcZRtDQ9ozcffJ11WmO
s8mqLcVCxfDjwmTkykonMw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9856 )
`pragma protect data_block
bhiyMUiNF5NmepQSEMjx+PAbldhebZgiHZeFONMTmn+bqG4MN6EMfsF5BG9tqKMx
UjY03QqMU6jgWBYy0doshLuI2kcSitOvsQbqyCu4mGnIMinKl7EhRXjQrtP4FVt3
F3a7ncAvQzEtZj9gmGawdgfYQyvtwSDmPdyIyPIZcpSJZ/HrdoH/ChV72THMPpVt
WfPPZiBO7/TC2PGFDbQ14L1fHyPdaLPFt4l1MjggydDInXOE2lsKgwbHuPi7f3mQ
SujfGa0PTFYae1jDptRuS6LH+QoYhGbhPcNXjuEeJ1kqEKXYi3KvFKZgWdOI0o93
kpZsN+diN9OPEEzXzhyz0ZVd/GVHn3aMphXgeNsR5IXNSY2bt4M8rns1UxiHvp1I
ZitO8Y5OCeLDanWRo1Z8M5TzTE/pkKqI7wIZKK1qIrB51oGKrnxaBwguHZDTNSc1
TV0rpCUNLie8pRncIyAHEUqcSkUC9bF5demXUk0VRNiDWoLBQYeRX0IrHvkZ2jEB
gwn9fGzheb55JXFZ235IQ9EeE6sHK4QQy4Opvy5xLlaeisPfEOkdhA9bEYu/E7Cm
wHeixHIoEVEdQwU1inlbG8rOwCooQqyIbvcw25QLY+TPwATfFZVx+RC/kZNDUyzn
2f82hWAJQ3xB8pcfAEmqUhkTxJhBbfiHLKYUlhoeeKR3BcjAtbXuzb4yGdHBXYBt
5WPIPxpchE0s1ADCPayhJCI6WGiStFKTbl3Euyg0iv5P+1dQUTQOPyPKuHjVII58
AZSV2m4L3rZDIYlF1omc66RG7WsCWdgNxH2Zk4o79WsD/PUwS8bmGu1BMyUVnD+o
llp29dPm0lnsWUdyTZ2sXnXypHTwGFPWMspg2O0wY5sKpsjcTSCnlveSR43OGtUy
yvY5sH2CToLdEjg+FY2XRU0aJkihgJ0hqPwawJRfw6XsKV6RaVyHDaULlahXmQGc
Mo0RZ5ua4GJCzifDRgacNmmZYlJo/vGvYbp4ATbq78L8DF9Ykz8gLmO88wBFlF6J
2PM+aejeifv05NBKnJkx4QhMFmgzEuxAZNadCb8gp9m/ngsRNNHBsw29in7OEzux
olrEAZnlA1OT1EswEutXKMc5sS592nPDLgAMcQcaJ/rSMvQFih3SpF+NmG4HQAi+
l2ribMzTvm0tC2E04gtLZIVhQkzczxvUzxxxscwKqr0+7N8visfbmDGFfRXMAWvD
d/XKIGwGVbtQtRBIZ95ZdB5Z1AUDwyDPpBH6j6P5PnptezgyNeQfitJNXctj0fE/
dYlIiHTHC2y/rLVe7Ppn6RwtiZpNGPXGjv7hZ51nVtRVNYdVvTOJs70vobtr2NY9
933Av7h01xj04Mmi80gRTgAejfWmKy/VzH+aZPPC536VgHIMfhBpzIPXi8Gug2Ce
6UQF1IvPFyVUjuhYRIw4xo4KKxTLC5ysG/C2JfjAR/7swlnFFuDPMkfCnujFkWJs
uVZGImb6u2RG25wScd1+SBBmQuB5iqfMhDb3a6sg/MIVGbAxLTnFC5BvjUb5IsSl
i7Edy1Tv2UO7tJvFLG6BM/zNKF1BNjpZ652VW8vGLDIHbMoNo6OcwXcW2frWTwov
oBCWWFjXvBNorRrV7Qwr6PHUIkBZw256z72ms4wEtVChKZI8yTr3TfVMpqHAaqwQ
bAorMWQ06GeMJtQnryw1c64XikDUHCAKh/p25Zj83Hwq6f/uT1Olch4p/FY9I4h0
6EzMGqFEmJqXb6BQJkfKer6aogjVUl2afgAVvhjyGiktrmhf70b8/7i/96fV3jW6
JcsMog8wpDr/AhDpNojFQVnj2PHGCA4TqlPcNNioDRoAkD6k06+yTubhJJOWS3hP
KUSTai+1xhp0Nd3a5yPPfFO2i42SwDwMOLiReo8sqIf10aZtEj3sMALHjF0zRfsX
+nWx/S1qDVULplfvvOFfJOn4MBv2e6dxrzFB7NWE3uu8O5EZNYr6wYYhMBexfUuT
9RZ5E1IZ7+B10IPgU+/Sudnp3YXF4UpxY2l1RflZWHhyunbjREJvB87025KNuh1y
sPHE3Wnldj+ksd13se2iePNoRg+FdpXeg7OGszeFjPqWNQH81pBENSsq7J79O34e
kbqdjXH4JyXEhAEQr4F8BnBYN4hqZxPW94wUeKa2vK07mjRtZh2nThGGcNX2NUYd
L81jgxZSQvRCaZSxfPfZXpHX0OBKaFNES5BFeLPuLhyaG36qYi+i9/9VBrbp8MYW
JmnK2MLPN1oWO35UNO4u6ZwwP0Y1RdrGDwXpIzon2G0ILaji52lQrFCTsZXAdV9w
pt4+m14el3hd87GMl+nYZ/2dZxDrflFMYhvYpDCXc5d7/36x4CNfBeCjadb3dzFM
2Os8tkozMJrKTaWW66k/IIcK+t82+mTWOnx/9znCQW5m2WrW8OF95nGeG5K0qjM+
Edp6F61bcrweuDn/EDfsH5k0wXJxlz09dwhQMz2UhCt41YKktrykMVFS6GnUmDej
CFMkO03M5WOe5YTYw0VEKKP+Zf8j4PYiP8a0glSch4Whxv9I00Shw/bpDmvDikcz
H+84O2a2rrxrGG9xUY72hWeeeXRuLivDAt1wphJP+37E2IRJ2Gzo7h4Ww+exDBSB
idpfve1SSOJij7pfLYSQIXr0u/fnvqpkXl521ZXuy1wRHcWSJwHn4x5IxGH/z9dN
uO/IML0ycRmKPll4YOE0SLxV3Q7cRivDDSxGpooV7W5+qrCdDjMkavyILG2cda7v
i8W4wzAwz+HAL6n2rl1LnCcfpm2c/PuN2kImdFhbU3SrV2zb3fyEIjqqg3zoJIBD
vZcwcDsDJyrdotxY10AJ9Hbwgc5KjZVvwd59ZcImnQd8xG0WZNEsuKXGT0jQo8HJ
KwiDVedxXDoNUBKAL6T8az5yh5NNjQ+8uFyzTi5OFNKMvAeT9IFb1yBiQhEA0P8I
4h5sTLrIXZD43omM+scto8eEumHayvfwTulk0IWiGfGQDgAGnpn83wwPRkjrw8+w
BxR26mOcBLFlyg1l5RDaeVJcFW5iq3FV20bv+9xw3GqIY/piP0t8/baYh+ChBrb5
HpGarPhTrT9/CBbLnrJCcILfsfbyI8f4gdVeaRKadl0IiZvpHa4ZBtVBCE4Bn0x+
bziHoGW/blAn7qEr/nypVstiGLWIkuCxSLpX44S4VwCDuE9YoJohq6ebSSU00otA
cIyc7eMKVhfAkXfKMKaEtVtiADcxoX3d1wjIJXZgM3j4QBA3V4RM6NRkMvZnuKdy
/BYaxuZmiv6IgLTCfjPe51/L+mgIi1NrCI+tj8EqLXP9PZn9VCoj8lxXmfLxBOZ8
3QvNBwDSZioXN8vmb0kE568IUrevSomJUFbZcG07wqqEHEO6LEFz1CdcaKEI/uVn
85b4NTom7hjUtEr2ewJa/MMmJICmxqEJuax0xdO2b9OEjdOy0d9ujhuAlZZ+uY6O
92hUf899Fdt7ZIEECiG6re8kivL0ErsUrwvmbw2BgDhtkKdcM4uVV7PW3rQj+JyJ
CpJr+yMuWZMQJKrkmWLsLUZCfDjJ3AN0VgJBup6bF3gU/cbwyttxsizrqrs+X1ol
yi3iu4Khigc8Sayk/7vP/E/YciNq9iBZI4GWwYrEUKBDmMeNo/k1MN0Jp1oY2BfQ
hDC2VZUMSIGud2p6t3rdAvppwPZd8JYf6SwRCTAMrDFI3837wc6n140IjWRERv4s
ZhIjFa+ZANKDexacWAS1HG1KOFr79iV0qiHG5O1fEDkifR5G/CDCfu14VQTjeq46
ShlRon2nSlFkP8fCrPjX9A/enHsYlneod+gWKvYs7w9OUCvc96LXxRybxeyhg9qI
xANSdE+KAZTwgSGRUSBJkFE5wU6yIXMErK9K2LKA2huPCVrI7k6Nn3ETYLbYyx4X
7y4Os6DjZSRUQOIcM2S78hEoOmCZ0coeUSojGPBne8/efgoej7zKLNzHGPYD+ita
2VHdSFk5OrlwdhZIkZeJQTiHjsZY16Wrc7ym2C8vOhUS/Amti5dgZj8UCHotHknG
ckzXFKr5D+GjKHprid7Jp2aDIvkI3cnTkNHkHrCLBeCUznUykfGloLJ/PwgTheFm
qmViSOtHAY9WCAAWabchhstIJXMli8MGBrmJpPo3VWxCu4Qn1aUmXaHSCOicjlZv
ByIEFHRB1ZwatzjE+4AYNuY5uMdTlAT/Jg/p5ideGJhybboh5LG0jLZUa3XrYTMj
SDRuG/BKgkkP+Cdgg6B5/27oXcux6YPzyYtjnExTD8cM+I7PH9RHBq+mRyLnCM9w
qzFzyBKPZiG5zbrb1nw5uTW1zcd37/Q6f8Xhc5O1k9zpyMQeQBthgeMGtSlw41Dl
sIsfR5Y03/EbBFOBrmpATL3tZkIb6qlY7ZkaOvNXGB56hHuT+gIlzAusdnf/CpRs
JS6NCh3+/JLndinfZmbC5nKjWRMC8xv/AMyzfW5yXrrvKQjHjIVgkT4T5KZkfeAJ
sVqm3aP06ep8ibP/H1+OLUNHQCSepbl4ukcmV2MxWwIsZ7t6Us5WFwhUoLruHevf
CdbNFVz1b24bnxRLmWjHW4QLJQewj+Tqtonj4zTUoDF83YLg05VXT+DsCVi2TbI1
98A3iizfqMhBcpnTHLkMca85v3xyqW92b2+dboQX1Qfh4+oX7gc1yeyjcu3j+uqC
haA1Fp1+IxTmTKojElZjw4R0uYSV7V6+fBdwLgOJYZRRDssfoKN2HMBvjNEB5sQi
71RHloFFTa6gM8SAtuFaGqoHH66W5eyRRkl0LjZJlgsbRTRf5KlToaDKuwKc5bfZ
gwR17CJ8KfkS+cPLhFqgK1NP+3acoPQDkap94VBx6LiuFL3kpF9P5OSVWUtdL9qq
uHD/YG/7woOM8Nv58RISkLEg/QE+/MFIwvkCZmFjKOSRf8NMJeotPk0iuRiG3EQ0
01ZXbQcWnu1EjorHXLK/GOBBVOHPH/sxsqp241R4qRmUqRKQhk3i9GhGpqgZVuW2
Dci//iNbql4DRvljZB6Df3nELQYYnZGtzj98ijzOQxees2pIEygnqfN3MtWc47mp
M7TfoXwOzmWi527uooHkea6gQX3EB7Obw41MjwR3VIpsytAGa3NGcQPVmoZ2yWG4
9RqO6Fqsw2juUwL4W3eGb37WV5ky+Lo+WwV6EiBrOoGTgHt3zEnAE4RIh6Um8WX/
yXyd/h3YrgxOA/QqPGRu6YbMtYZswC5L/0+ZDkZ8bn4yPIlXhNM7pOPnfLvQ06+Z
CojBl+SqRb0kYeA5YmBWV0DZDl/6xNW4tc4sx7FKKbhsQxt6IC4OA3dNqwhO5f0n
XttONA4rRrkudeWEVG1LIZ489X2yEv5BV2h+Cz4dgYBRQ6i9PzU/qddi23rOfSDX
wbKNRkg2Udw+iDW3mjiBPnckyV1/D4a1+P2Y68QoXlSOhuzvKxG+5WfHd+yymcq3
zcoLhgXHR8NrZcfd5WVR6r9iXvi87XoGLVjtrY4NEYBB+u4Mvx/JnRBwJrQ9y8tJ
QoXuzTFzlB8J1ZvoHwgeiTLfrWd1wlbunceZXXBzSAnpa56McnyXuP9zU7vL5G/5
MzryqK8qTs7wKdRWaewr+G8LlylfEk8xFWV57Aa8qgY1+3Zx62hitynhSPLgDgkD
8JWgtJEzf5q40XqECV3qEQJ6pa3+aO6AEgOCpI/EVSqKsyE/Vf0oZvDb3Gpw5QQQ
W0jBEzaBFp5Z4+R0DpF6U4mq8o041+BbdA/iDz125wCZaH2/M7CtsMrwxmjJDa0d
m1VMDko5dc5hWBGF/7lrwHRKIhLfWckNc5Izg7DhbQAvaET4EDOC0FqLQWnYiGcH
UOume4FQJpR51gykBJIkqhVT+jdXyjZlb6gHXufWA4zZLxIxV3IAQCW+mSudRxeF
XayYDEwoBxujVmtaFtHf24wmHtTVdTwLnVodz8PoI82A5DT556nSG6ZbfdtCdae6
t/ptV/gN6w2n+5EGuhi+BiXC9Xco+kWFIArmXERxP5501yUO9/3qDP+MCOWEpR0r
M4XXRfcX2SexycOXIfTcnNi5ZPqHgyfbUpKewrp7+GncZ8xUjNr0zOv6E7XWE+aJ
A9GX6ysQYkrtrTIvl2QdZDaEC3bUl2tkA4wFgtw4EKeLWlyg+sr60e+GVwtzjKXT
5F1IWcqI4L/P9adsJgWQ4s8zE6o6U0wChBbDYCH/ib1Wg4ysK1jRMRmvB3P+HRZk
41F9J6BHcItqlKPNmhcWzY2VtS2CFgcvr3JyVAoR8wmE+F5vbBrmjZt216BJzSf1
SSbtfWUy5q4+6Ha9E+AnYlsy4QZ3fSc4VWI1dNIv27FWUFL1BqfV1I6wB9hn7CZR
i5nYh1MoH/nT7xn/mYj2hHriUgNhGK9I2SJohyWLweQeJ8uVhiZJDEXRJRet1QHm
hYnYj1zm993ElfVqqBi2ujNqWxd3BG9n9C5a+yKtjCDzXqwisASn+ej5QRPuTW8c
aRCKIf88FgKeq8bA8MCdi2d8ZzEwkbfWHcAX1FFmagW+PlDTuec1wISR0ZbsDz5J
FPRrkiLRSsHMG6upHnTwCTsdqEthFCmFMvupS2tjQKnvB4OqzWTplUatgbujFiR7
4WPp2ruEdazY5ne0S/UBsN3Z+NpJJnCtqo6l1jCmk8rlGbGDs07s37oVfCFVRSUH
Ox57OXJLpWaiRYcMACjZpuDiMmVKN10du6YWRb60B80xpN8LWHIMPuNdDonx9sIg
AF8Ggabr4fRTw4htOoNsOMK7pykyKLjZWiBPYTp2lJctE9viKtJX1OTaU7bxsRKR
YwXwhZBuw4kVwS0OoIXceqSxJoN+mYoGD5g7dW4G+te2hskuS7ykJg6OXD8wXjUU
VnRwXe3ao42F7kIhsURRTNRUwekhsz2djs39iLxd7QFtysXRzwfS/Ttm1EJTwfvU
4yrZgT5gDCmfYVHPBgubqSFdj5F641mkjYyZMzsrPAiU+1mFXTpUhcVuJSghJP7b
A0IfWJJfP62FoJBvjB1j83adjt+o4YrlFNDSGtVaVtN1Fz2Z1L+6pmr++juNlFNu
W42ozRLh5sCVNJxf+j2r5oOU1eVImHRBc/44JezRLaXpzcxFT+9TRE1139OpQqYz
hHehiUgrfGsv+1Zmhao1q+CQ1BxSNR3dP6MhEFT/3D9NjNSxVmZkb5nxQpK6nPZL
9D1ct/wVHhCuPEEt/gzSJzZICRXzjRcImCEzUdMfwyPdV6AN0HUlAsSk0oTi39il
h52dHIZhGGI5y2HCUx2HEPfIs7iq9LqWfqRYdKtBsxMg/PUYoifNKGIU2DzuIYgB
fQM42ys/fpFGNd0xhU8JgOxadtp0nsgRxNGHnF9ZctixpBYC1FsTgnfrgbF8Xis9
eBagATNIREFEldUJWsftJ2FteaYbniTPecjUN+S3hsEkjYZ0JrvTLgL0lLDbZJ17
GJ4FlsfJDelDj/HzhwlA2khSF6/Nx6gXQm2W4Fqf6DitwhNt0ZfGKiVLxKWQ1rHf
r2RwAlUtrzxygKKVna23uIGUd5qRJxYnBUUApQGUGd7E8qwhchCWRXeFv/1MB1jS
fMbxtpQsRC7FcOWbZ6sJBQ1YwgebyFSFg2WPkqcOjLyl0ddDZJs2bkVQJ4bqR7su
Rul5+DpDTRzp5mNHERm/m2FbWgTDWofta1EJVXCIKcVNDlCcs0YyIILd2uLKrVgN
Yl5DszgGVg5d+W8dIaQaEFkPLXU76vCH3pF4f7OhkISjTmigl027qFdyqY9M0zGm
kTvLjabuzSDOtcLDyOsPdVuPvoY8TVH8Eb3N8BjSdWjcA1PwfKTolzhRvT66Y6wK
1MstymLlgHaG48br+3VytDXP1PcrJ8VSA8VvGy1iz/eX4uP6109BmX0VGsNG7w67
LuJ6xNWaUGZT6znhQRZeeNcJv/xBByRiw9aN41K6mvTYhGo1oaZqs/GHm7Lp0lRr
8dbgmQ1gZSWguRMMlkMPLSY0lolD/Nk3/OCgK4xGnIjCizD8KP2kiBAaUqGsQL4v
1XBWETv9LoVWX527KNXno7SAl2OB8WfSWBzeYMqGNbanoFLs4Fs5sKBv8laWX0mW
KT4IuSpS+Rj2bHrLP/lgvdVr/ymC4gIBhFaoJbOMHBYQwXqDxIN1TQ1QK3QozwvP
5/+34fuLe+m7C4Pj/WpSDQC7/k8L/UXhmkuAEexgOqCiLH0Dojc0mOBJ59nTFqEe
/NKdbPlEyRr8zLKSThAMzluFmKm/YPVIKdU7pVXuLCtRAGcXAxhxTlnJdiVV4JBA
Nu5eAMONzW9uTV4jWYrpyv3NcbJP6KmdpyziMbURuGLVpxbOD4xbkll3N/S7J7rJ
6HcFX9+YXlZjFUdXmT/HoJnb9mtODqAzldwxFbuB5CW/umwORHMN7Zq+jZ0qdlQV
FtEiJZN3G7WFUfWfLF9xqCcI30MLsTN9Y+FIauw7+VKlzUT7/VeDl+JFg0iyF60F
2yj1ldSJ22HqSHxFZnN1hmFjJ2yaMTgq1o2sFK5BNGRGeiIis0/7SrYJJhDCkmxu
S7ckbLtVIX7kMuWSUC1THfY79XvQ8WhLeGMIR+nzWu+xCtEWHtKbBfmhV0mFvut4
mMeAwDAlYf+bgrjwwE+WXZW412iBdEc6merOiyHYn+I81ZXmsKqIYFt+NTFwaRTA
FQOwgYmu6TWbe+t+iZWY0JTbrxJbrvkb1MqwyFWII63WfRiekG7apPx8XQOjSDFm
CVwZdcmtSjRZ9JmQ6wT3CDJu5aAkWEFeb+2JmfvBh6Dgd98TPrcBE2hEMwIpZLX1
o7WdlqtYU3nY4vF/9yKbXiUq8zuofaY7s2isxva5AZ2Qzdd1FLD2KUjUFaq1MNXL
+QgozvZeVVZocIj50B4dyF4cndUWa9/ATU8sYsN78w20iBioURml7mhaC9c4N8m7
jqdYQen7lTFFZxdlihYMLkYJ1zbpw0c+Euyf/3TXe01nDVYbBFfnTZe2aVQhIWGC
toXtLvxddyOuigvO16miBn4AVaJ4EfmMSPz5witd05otVi+7QcMfSHxyymlzO9hB
Eb09Z2mF2lmpgqs45upRAnYcxNtVM3n4XhwgWbuMHPSwKel9rb86NKMYjc0a/e34
gDndHipv+4fYJuH+z97HGf/6NR2Y+nr1IW3kWKRAK0jOj2jJuTF/p16gMfdi5pQI
xT10B4U9DMucBlECsbzCfnnJBQD/yCit/HY6VHrKSC9+VKZWH/cZYkbaP70k6Ovm
af37Y19mudaKnMH36TDRmI8Fr1bJBuFp+qOXIoieFvRavlBcKi1rGAJ3W1Y3IJGT
X74GkZohFuqsRb3RzyWE+MSkHlCBrcLhD114D6GH9am5cmRChwYIi/Xp8SMJYojE
kGtQteDowvhAfGjlxFd80UCR9RZWlU7exHYM4XtR9DXChzIcPeKoPH8JuWDGjdQ9
j+mlnqyPb6SVFeeUXWN5zqXqIi/AkcC5OFRDJ9ysfpzStvsw1g8q52kb6iUzaNJv
kqON/hE1ipfeCUFHrUqnzYo5+vZLqcdMqGQbvZJujdFPOr99xsCD93DkUUUAT/13
wBqZJM9aOhS3j/o8NI2aPBdYVJqyz9a8PG4a1BJi/xASZ3+opZXr/kD7qly2Msa/
TvXMHSJm5Z73N95q8BXB0z8iYeLPEgmfDi2uB9k4kWC0o9CMqklCvIsp4l5OOvFO
TBJD7X97WvGOarpS/I6hWDZ+GudOwK6QhlpiG1pBEGmvn0JRWGQsUzcgjMoZmruq
gcegOQ882SKPYSR+9dbxKd1hAuczZJnR0/SwEOwBCE/VzRAhk4cVlB1NC9D1sqC4
kTodOkij9+TW7m9bCUGSp+pWiPV5nK1VWVfC5m4NHjEixzHV54k1DuJM52XVcbW9
M+bUFxIehOzXtCuf3xQoyfRgFCvc7z43IOFUGDOlF20OMIYVDtyyjdL1rPSLFIPz
NVFvayrTlBrbJsg0ksijtOIeEH+5Xa2C61nMWKSBCA9Ir3q0parYBN/W6d6+YJF3
8d4oamob8ULS1eycJh7prG4xHdYGI9lAUMHTpigVnc5kXCEE3hQik47xmxYQAWFG
fsF54bDqJ8PiF/N4RLUkU0yTHc5Ixy7nQ2Rq1vRCX9V61S0OACkvOB9iRd/ZFxUN
V5bew8hSQAU9dItPegihbku4VaD1BwgcuOvF7yVYanMq2xqH74Tsha5XA3OWntBS
MeDDLnJz9C53B2G+mPry/RsRezPwSKFxzC6LAF1SPiOj7m2hTxqAyT65TC0E9YKw
GEBAs3AIF9Ml1AFgkGIbqjgOyB/S3FEzkWZ71u6StJ6MuqN8PRUghNLEquKB4GdU
PqGjwpn3RD6NfhNKnX1d+oQAE0+OWsJtpyceRPDtXyk5ciU0ToeXW8+SkNvkAp5O
O3EdGYrJxBNZeqi15x+0+OU3KYK6ikNKJ1nS6VVVw+usHbyYLfJdwFc6jnqYfFK8
t1MW66ZnE3kvGkx16/+FEJDBXB9CV8/92MLiKZtgi3a6KMYXfc7qh/TMXbUOn+/W
pKuhLVKkTB8o9XDj6EsY8rGaEALCl5Hbn9jO3VpbVruLjV+5qEswPvAgMGbV0rwf
SQuEBtMcIHdFtQLEdTEjCHS2D7Y+6cA87TLX9+QAkY7tMaX7by4g8BCb4XX+aJxB
XJFVGKG2JSSGyqh8p8bDx0hPE12ef1ZavlAeGuuqChAQG0cNb93uu+403oeBotxn
v/sf5s6FDDrjaQXOB1l01oOU/ZsAfWfqnVrAAb5lYDLkf+mnmg3594UsWUh/TxCC
wYtZqHJxL3CfqoWDG2JLI1jI5Y4lYvsG8xUbUQvdKVsdAuCiD1INWUJ3prOVALgR
JG52EWPlK1sCk+L9e+fpJc1VlSUdPuHHkANIDfCqL2zHXsB1aKRBqKkDmAC4IO2d
oeclJqw7in2ghT8Bqc0ONWi6OtPWi68EmcP6sAUSIqkXzwDPIkWOrVqtroplR5WA
NJOMnlYE4SDB2Dycb+BcooFuSXaQGKPS8lI8QMpujGcs7ZfFJgtBm2YYRM3UoxXn
zj1S6tPoYTfxrG+N7z32poD+82IHNdLYBORGrMEE59ulbJaxhv8kf+KdY3y6C1v5
EkQdHfG1rGZywvbz1ER3WOr5eEvWp/CixYIif0HY4wwoloXaKatcdjwepIg0VKCk
vz4jgjqc2sqm3dCYk2OE0BrQ0u5HwNsbRvGP9bwrF5Xr/hwj0nNEnzHE1alwJAkc
s8wmdkJ9L+cRIHKBpmQXe2f3c0qBaG+RRpYQRnNZXL1bxEjX6ZB07nzcHEQi3NIx
XnhS7MpdN6/xOm1VBM5/YL20y74DNamuWLdIL27coLwKlyvydfbH2yWs1Ls1u7xe
G240WnctGbH+NTBRaulqGg7HVuYopKFaJI86kmpNFlYiUj6Xt+YgvLU7913lBePU
/QPUqv8reoLgrqN0REN822bZXngM5MIzwb0e1dS1pq0VTh6ENoLfDzHuyX8ONH58
7eENTawKhK/GdahjxL4oKV7osv3XEFKWR4U601vCfWtroeVYO03zmxVJ5Eg0PBoW
p3A/B7DR0DlXVUEUrVLJTe/vY8k5B2ol6jslvSQonGgAMXCpsLu6pOJCInyZESsC
JWOc5Ht+dKYfE6w/659PRbxY3vZ6IHg6A1PFG18Sa6wk+ebLJY22EhRTCTFodjHb
ezBLqHM1trpk+9PoLL4J8+N41VCcsvGusdhiR+ZUAuvCZ+pMc/N2yBR7Mk5h/Tey
5rnb3UkRRqtwVNukTaS3K2FTJAiWqrI6gyDxilUKV3VIFLD5L9JpfSmbwui0wQeE
RFNo2LZclbEEkxgKAs/aAUB1DpgIPHFUDEZSJUlcorjkO2go3VD9sz2qxo8aLANU
J3ZRyJuYutED2xkfVtwwSgaBGBNrMiqorZX8sz0IlJgLnWvnSpLr1Visko7E5nrP
2kHyrtrbhaWEtIMS0i268sKZShy/m0V4nVz+pET8FzSdtT4M7n+wGpK44ZIxJoXI
DVAvMqYCRfqCD5Cf7aDGHK6QpqNXKlKb1xs+Tg1CMY9ZJ9r8/PWkFVrY7/pLCNlZ
bV48xvAyXQiftu8tTUUAuHuQLwp+VStGb8PAzWPWUBe7WTHloRiyb9dBF+HTGSl6
vRPuY/jxZlOH9dqLN9el+8gh4PjKmB8rU9fOF3S4SAPzmIioxyftQE2MciBPZDng
rSdDBdrTyQ0qJVyIK0ydQ9F22tzqEJQeYCbCmNpQq9VhvGfu0SYx5Fu1ToH61ai1
sCsIubFr4bRmacLzbxwJc7DGfE/y8WwjuWRBTJq9hVzdhD3eGmCPQoN0Wo1SbHte
Mj9xRDtDpuwQaubjMwKrFE5tiCu8creJx9hH1MUdKS3szEbPPYwXQjawFhhIqF4Y
XxyFxcBwCl4dryTLqkICWT38BPN7ERYE1OoSEpCLiFpXIWhLxCXxWqKUajlfGaJ2
MOXRcKXcAuRdg9OL2sZqfzs5UttbsYNMKmw/KGaauTxZ3fvDPC0GBft18duradL2
EKnLK3xG21s1+eduJ42OVnr3SQ9sGIqVSZN7j1FL9MoCFM5PzgQi0KP0p701QdDG
3NnyHEhC/ZpKv+LT5wJfL9r+6MGX/NUXDlZAVJG5KJjCoul+sxgY89GiXurKNszk
sDwdf9qu0+g125MIl9GJntS46h+/k/GMKNSlPzit1NX5kgwrFLsySTe58578epRb
YbCgvhr7gij5Oa0saZxTRUD1cOGaOV1rfBElVbIWKlaBBTn0YartcO0AoL9xzTJ0
UtkDFW+L0pB0nWd+Ci1aZt8Fr8M6KZsYVl5BciLx0wEfrw1/4QdWp91AbboC0k4F
dRNLjeqkeez5WXpSti1cSfnB3sClW6yi/XDiYQ+ESFzGucEHkiy4f++InE51Et4S
5dHx/mPBut6CS/fZEQZlli2fwzWZx0WNTj2UPKTmNUi22OHs1M0dNC+rpkXQy6c1
YnIwzEUQuyU+lhTcheIXvmVNNPiv29GhhM/VCRcrXM1CIlgH01jpJZXBIeRBvvaW
eDAGAy3QF2hr07HV/n/FwLcApGrOn+toksyeSL5ARIJ29v2MjbKt8dEuHMkGn5rS
DWwfp9fnuSD8EdYXZkB/vS5wzAvATcBfvVEahRMqlbdL6cmW3AlmnrDkYhOAaJxm
gwzvcH1Qp3uCa3/QrVrlzg==
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XoQT1YCaParkWb8E8bZjjGX1QAFWjOeYhxNgIlvlka+yvmXUPA0txgvquvrKjsfS
nsNR/w4okffDuqsq5o1SSIuxMW8ipsLXtUTlkxHBc+HrWB2xqpj6bu/LcfRLWOqE
voZTREqILH82SyUn+5SOcMvX1J6VHmrIWO4aaeNK9LE0QANi/60/wO1gNmXQ1oMn
nhZPe0sYVKFjjfEh3PCSf8tR/cm5h+AezGwTWxhOb647Hj4Z+bCjNgDuRO/AAkXe
QWKYUCvBto4DE18GYngUbMFqZf4vRuWMU5LXXHRnT6EXuSi9hd3x2PvcZ/QYITLM
XDObKzdOlxPsL5Kyl3Y/dg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 656 )
`pragma protect data_block
lZsK+lC4x2ObDtI26J4rMbtrk/mh6aw/GW9WfyCZsbBaMSfuw08VN5+0tsR4n6Zf
SX8VevfMqiEkHEV0ltRynZMtDD5n6U4dZ704lIFdMQGnJ/zqlyNb1ujdch4RiEof
8isp8Dt8WgtaUoI/6uni1eUM7IsrXJEMviKpI75NVH8j18vYrGGNO5Do0EtFJkgd
j2OQ/dk+qjwjNAA7i+J4/pRHhOAdtW4g7MCDnXymu5RdT8wlQcDEs4OIWUH9Q/6w
DLyLszNtbhjK9MNssKejEdcMMofs8eOi0RwlcZVYSKizQ745TJwXsnsSO9CKFgPA
tIo5GKkAbKVW4AfdYgshM5ft5AFSAa+8kNICOGLnHCbWOubPQvtVdMDhE48oih5F
ZXSQrGB185H83B1QZYWc9sJcL9GcBS6bRvsihms23lvAmu/2JHvSj4d8bB2HDe8Q
/Vg09X9AtP11el8sHwGl/lfOJz55lrvjTpb09jBGWaITZMKee0xFmjbqdpRAw+mN
TjrAMmVjNEIkCRgx5b/QWuNKor0G3uB4jvZ30GeMKSc6lSS12SEflOV8LumqJkUh
X4a8ePkMcXNTo05WMNMrsUjPZRu4mD3/Uzw2/j7Xsx7USCQPxjlT6G5lByk/AKNo
H0iqSJkP82VIYJ8LHO6fp3I9YznJInKTYM/OuNfWehiAZJoWYxWmQ/h0h68f55dY
bcwpSRcPE/rq7G3VUtXgUeeWrAfAml0hXb9LmLjBvaVZOamPOGXf/5KAbhsMAAqd
9Bx1/a33uPPK1NIZBTymBFJ/1n2uMTCHAUXncHMytKwrxk0/WHYMJnar2XWvWDWS
m5BvUqsyMXR1dtXHfM9HoHwgTkvgv6mVX37stbd+fBo=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Nv4BixcN04pwVa+/7bPNUVjLvApyvImqRYsAONZwKZIEc2drrXkukS56cocBP/pM
glZEEItAhcUw3KQWUXbbzrB+RNT60ZaEATObPc2FYfGWTWF4LURSvK2gGHoFfry0
lnP/Hz0YIV06hUgsokvsogLwL5aOA5svgTEtffLNEEfRIjV6tctl8Sk294hhpI0e
ruQ2anHgj1kPPEqpeudvrj6UUjGS7JikNUxlZYwpfwPufLbF6k853cJh4lcY2IXi
gCzEMAY5A1clNbTVPLyJIRIr0JXf72dP7kzIpB0f2sO8z1GfQXA1WhiBKblTci2V
kwvUU0E0FxPcxlBSE5AGtw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 13232 )
`pragma protect data_block
TtpmBGnHj+uKET2DXUSe3+RgvGICIqDc/pxqlLljTEMT1Bj9U60dCyDZqXS7ydYq
/tKYQcE9Amgu+XPajvguMIOEeER3vkfsjugKqgRodH/fUJsUnXmzNs2cZzybb4//
3uqy2W5WQ0aeerfBJsu8bRuJPZ7/PJTAPvU0LcJFwxtWIxCOhP2rpn/XuDIi+d6i
RqNEh27oeiOPR+dqA5dLnEWVJCzt4MYHNSF96HSJM/ZFL1hwSPGLIlybwwpcq5aJ
ziTXTzZrqykIm57EgNTIV9mSUgL8EpTA34QMwXr493QrTAT8kQoRv1nrSaaFUpcH
S3qzf1MRBWg8sjViLN5BnLmzcWFjuQF6BzpDM1tERksv637n8S5TwHHLBp43oKHy
rclBmdGi13Uo3xss3FbEKSKKbWVRCJvDm39TPBXXT9vQ+FDN1xqsmZGojwW8NX+y
5BqkJD12CO/6d1TDwEkbkr7o1H0Ow8dDlgAmsVaGuXXb8LsmZXOthEdttyRNCrKp
JUVQAwBaD5KR7/JuuEp8iYkH8uEPk7zlJNWDeswz/wCv3vb/I4+/BAdrLf7S0paY
l99c49Ax7s01JsAXxyI8JOc4grNNmzAM+jELGDVFc5rvVNVj5wgB+uRLtWi1g6cn
B7Ix5UteX8lcnTpd2/tdLLDXUM+qSd80F42VnroEydohfOUNs0CU6gQYZ0L3oUEi
XCIzapnK6mG5BKFIyyp73PHnDtRdTmm2b+27CX9tSMm/68BSY9IWDMqwv8j9Fs2m
8cqj37uxklR+2N5pRylqJyf0s+drv7NgbX7f0ISD9ngHj3yfhfMZ98ivFEX2gD4j
YMT/IS3u8zFKM6aXFGR/fpaZ67oaz6eVv2FOWPSEAaMDr1nqgMGVhoD693NOnI0A
bP+GRUX9lnGrfkf0qyXgFPLkE6oIRVijXjXUkVh7NcUsV/c10GLIFLWt/4yWBc9f
yI2RRNQbChO1vHUjgQeSjCc+KaXZ3S3720vaNMPHehguZQvBInlsRKzWvjGG6PX4
H9//7LR7toI6+f+jw1NgsgmhXTsnXWitFrSYtD583DS/MgCoVmjHA35h3kKQqf1X
S9C/YMVYsssnWqeHH8gDjtntmsom8uIBmIie6YjeoiGGkzSjRXkYy/6GHmAPNJ15
X/JrAc8mYn+vRY27CzgYfo9sWqRroAyPocrmJkM2v1uW1S4ua3VDt1mXCTLl/kOH
xZpOpqz75rqnAsHzreMJ5rqROXvSq195G5V+tMk4iJ0rUi8DVIhcRjmFB7i25Nba
buBwCicMw5FtZM2DW1359qWZyIiLZAmC+ESNA48zMAq4EP8qC12GieiFZ47cggrQ
Pt4qgeGcueDYeLYF/6HoA0vsbklEcflUIG+m5AbnbmYYzL6qCEAJmZu+0cSc5JuA
JRMcAAu5zOGWfeXvCTrrn/fXb1E9h8YN3wVkOuJC6bFwzZMII7dWjU1kMWc4jqUj
xtMAzxzUxLcZtzxMYGw50TGFiGcud472UxbI/LKxu5J2dmpOuAc5C9QeCcidXGe9
bgymLQ+KTt01SMJu5x7f65itpVF0hNlsSEN8AeBJXLK4sbyFGODKPQPHjPNDDtdZ
kzgGOPzxBbrwvX+BfqK1dwsrwSeadS2nDi6LuG02VMALKtdL1QVE1DoisVaLRTo6
K4Yu1Syq65dEHzmK6g5Lvt//4Xj4kwKcaPt2a2sD5Y5X1mM6CQyfoHLyiGnXUez+
IvlQ2zQROreXTP+6xkXp5FsdYmgGN51EQAWUqOkY5wBvH/CbuYwhRcxmq4OXO4rK
EjAJm7hHw6VrhUVNflwNu4jYiBIceNJ2dvKt5/KDFld5j7ejfjjpvrLhxfP4V0mX
b9FmdzOhnzIBGQVZUaG0FXI52673EH62QWHq7wXyoOY67b1SVz6mWegZZ1YgFmFU
dcuB74Kpar7yZo0C0GR7MYGOLsBEWYVVANY39KtEHG9qQdgFpzr67tLoyYoDEYfP
K4QjPg0OCPm7luZeQcXYlAiXVkMi5BhLIhGtjC5oti+Tlo7LEJnUpfbqf8wOHaXo
rMea2yI/8sC42/OLrTuuatMMSfwDsKosTMvR+sJVuDbjkAQ4X/44SV2lNBPDC393
R2MnI3X+4SyhaaH+rue/H9EXnnGDOHfFwHASbFE39EVJw5pcdzqidrFsBDq4WMBi
YR1Itle0yqnLb+qvPRcba1XSE+fJR0aSiXKmyq/Q2owjjV/Ps86ZOi/6oD0T7Q/R
NcuJCu63VBxsx/bnqegmtbEH47mNSM6qmFH8XBIBc0haS6ul1lvx6kbLafxZRXex
daTDpUCKHB93aEwgAnaYEO9moEgCkPczfwIbwZnv4Dnwcn9K5fNLnFZ9yASiMsTG
P7RECoFgFikNDrY6Wb+KVuER3map5bQPZWBXbMMEO0xtiNs8hWZRcv6sl+JG4aIf
aB16AsgyDESQKs/O7z8AsXrv1t/yxaOFDS71rVN1Xxq376tK/0zLd1zF3MKaIZb3
0cJwv938Ap8HTyGL+4cPFiSbUZheb3ovb5hfaENy4nRMby6KDr3XZR9cNnklh6f4
XfE9tTZIM0iJMvEUzp0NPyKm/4aaA6LKR1vK2zNDwhZwr2vfx0YguP3Lc3y54/jx
enbF27mJx/oRWTzeMew/61fUhl/SAkT9DD5Mtuonv/EdbVwYSETZRvktlPq0J6lq
+dl/0ZwKsDV2n+9NXCTMsGDUCGe/mfIk1i+pswt+5B7Lajeb7jDtKUeVFLvBO5de
iqXttDAw5aHENCpwB0/D50Ns9F3fIMkefGTxdT/hWHfP0hCoB7WvdQusu3rZMd5O
lzBWkGYEtcC0NMYo0LpqF1gZwp4kMJR4LTsYCU+xTmwYCOsh9gXWL3EakHFldc26
bb0B2vENX5QJJNfqIrLGjBBJ0kyLlq/6JFKWkSq/StfZpFtPUkexPVTHQHYibCBK
N+9PUGz1D14sTIeyH6u0hrcNm8n4cbAR25v3yaQMqkIUe8yscM8JOysIZ/1yhoH/
rNIRGA3D0Bfo7WKxdvThf+cewULS86kyYFus+GdeUxC6BpGJ6F4iyLJPJo/cyRNn
F0DbfqxGYf91sB10g3xX/EhOTn7L3bp3QhwNt8JLYmPps/kAE4R5bJlEGlis4P7R
bjvIGBhr7lW9pXxNxd575Ciwn0mWfPbY4ysIcdPKuPZElTGIC/i2mtJf74OvuMcj
sj+FFHcZ08hy/wEjp29/+r2Nei3YfY0vDYOUYwwhM2zMj45IWH32KWkdJY2Z8/5V
3t3t+ylXZ34lonKbmLsKxp/ILcm1YYu0XIJmpvA1DzBjo6FAL/yfQu25lp3i/EwZ
m7WAmV40q9Kq+Tm9eQMiI7lRF/GVvs6WBF7OIu2XxcntY+ikFGwvZTciH+kvgd13
S1KDH2rrJb/q/3rz8kFGFRJptTKlZPKRrmS5qh/fSJd5dq57h+DyDTVn9YEorRyV
oDuq+6Q8I6q7FAzEqmq0jlgJ6brYT9xWc7DC6MK9CBsHF+xlwgmrRfmn9MpjAy7I
9R6ofX3C1icSWqZVNQsVIAfzueIDLz9QRGkgGMCGujsmdA+k+WZBjp4j7UoW6NJH
5eVnB020ZBlfSRZtimbMjs3zUaSWcz8PyB0aHMVwNCtovfnT+5Hs82aJ3VisNGx+
6oBeUZR9jd6O9Y2YHndoeqLR4Yj5asE4JRikeCRVJFo12gtWeAVUVFCl8r73tJGV
RHR/jxXeYvTsr7aRxf+ne3Izw34xrgHJLSaezM6p0l+2xlY1T6uaXoCVO2rqMBT0
jbQhfX1JnyprdYU9rMFlvtjUMc4JDFBUkOuyTzQuLMr1m0oRS6lB2CdndTbzzuHg
0+LQgnbZP/g3ltSEB9o6wczz0gmhkupmXWSW5y9W7ROp176CJFuFAW+/j+yNzdhe
T0MKp12LjufMFiGBgGEwJWhu6RfPLqhMDEizWFGuuN5TpliC18DHXWdx3yhV7M8F
KlKJdUzs3U1BgRV7knbgSflAqe165kKng16+poNIdpPHmrw4BSAb/yo5njixP4GF
rHHEkyy46aidklr0SSLJJqKVyiFXuUAB5TuzE+XQZ1/zgccVXCW3jlnoQSw5TuN6
eHnRlkNu6HDJNt8PMJiQWSfrvwkFzKCSDUahXHZUjTk7M5sHpo4SdYxP/8FLHGG9
YHL4nhQLqUrjDRLQjJw7YtFwaji8foF3Z43mIP35tja9yysNq2JQCMjitu/vNWN3
51j53/9pHifqAEtdfs8TBWOrGjrfUoSTpUMMDR3SZNO5XTyLXyFkGRdin7Iqyp5K
OlDQo6uQ6rBORx7SnxeMpLzwq4+8x5VbvccR71y0hJ3IzibfUZJLU0eW0lrprokq
F8U4DMD06VSI6NR51ybBcpVKjIbIQTU4QD3aEQPiT6Xry8lMMyXrI0lgqvpAxnDb
Ep0/caeOiDDKGB+lImbNuVBbSlwRL3OgLz79T+VVrs9oScV6IqM2o5UtSHuzrmO2
WSM211TYA3c1xYPawONuGmgXTOdsuGMEouzIqpkM8yrS63I9N9DCCW7toO9T78Ug
Ft65exRxyeJLhhECi/Bt/P53FAkmvfQjlSt5lCNnGeSA1tpz/S8Wluazvbf2frAH
ZjX5QhtT2UNZwpLkfPeMxMyvxWAiE/DQ8jVHsgjXsVvStUVSWcC/Bt/U1tGh0qQT
MDQPQ3b+8AP2VpUaWhi0pJ+MwvIwMM0LdfuazzZN2CvOxh2OL5U9NV0/BdBRyO9L
hZIEYocZ2xTcIwXO+xAODRI28mnKwI62Kyi93fF3sWDsRqdS+Kmx4FS8mbckJhyK
JjPOerbz96nBp2bfOaerOQhyWk/TBdgyPowfNXJ0iQ6D/LGKeoDsMYa01xQAJ+x6
6gLbBC+KDrcynrBNzGPAvaURbQFV7NFaxKkZR9oAliWgyiC55FhTYWr8LJ6Z5Usg
Y751AvNfl0ViSY5kqKptIvxOenhIzxnxdMuejjmnhNZ66TxeRPKIXiOBFwvwiGy4
lDcc3Cxqi46OlDLdCm8q6wRqQ3TEHRkwMLZR/arzaUrbfCGP7177qTxSle8jM4i6
oNoEQT+CPPTbDC4xaVKJ5iOfp0h0xZq7ugJLg/pfWa7H4WRB0qFcNJzXBfBAxVYi
jfDyP47tXYXUOqR7fSqASvISTx2Y6ieOu0Nxgf85DH5EhJtiWi9Ng9dmgDlfbZYC
I71OpKDq5fN+fdisDOoWdZCU3JDtaxd1+SKFQONjewLagDwGo1HxP3lRAcsFAmni
Ga0Fvt5hp/Mpf2oeBBxtdNIedvKoz2Wft3whgyOCxAMR/VmTC5zIgUEcIh2iIZxK
/BAc0QIU8zDhgky938t8E8DdYSZuwrGHGxxFE2+vOTuKCqBuhaxDZsZQhGii0ij3
OqZ8nYrHQ+wXb5Lj2StbJTx/Hu2GucsFMgo07BaBOqvKI6T/2GUsDX5GZs/pBOj0
r42nVJvnqr+xTEyjM8J4slRBSE8sKVZZ95g8YxmugzhIwyVUDBxhGj2rm7ePI3NY
UtSJOaUaox7FPctblyeKfn8Y7iCLKL3TmvDqMRsvt1JeeEXFYWo/qNA3cqS7M5Zi
HojKNbWOks8ciYIZZ0KOcTryqYg6ZY7NhmWRNTLSuyIS5Ue4ryb4Nn3EQhYP+B2j
ETiVrJGS96iFB/h2yan4rM9X2bJYn8MsNcubwgC6CNWyYoIm6N8O76uKZqpzaJmh
MiQvA01p3eMRumW3cLvgm/ToJinagqU3n3QOQ4c7Jfzeh6zqa7NhjPYL1ZI85Dei
JZtI8MdVxNLhc1CA9dC015G4Flz39LMwug5Elt/oM8VGF0mExdjI7L3U1DRyh2Wm
PjWRdbkG7E881RflooEZzlNJxe9x732cdfrmlYtHQPIo2OH0wSqQcC9ybXFr/w+k
x/Pn4DRkIRG2cewkghRDPtf34PsYGZUp9AkqICU0wRYmgb8dZAo02xl8hFlmToWP
erOZFLeXqvcrUdsXbSy4OMh7fWE+DhMeLp9oig4CrgZGNq5neIXestVd2qmrX+oD
PePCfBl2YWi+XEW8ru645iPJFeho7Oe5l5T5atfOF99rPkDgWmCWdsUb7FryO9fJ
gqQY5vK9DkuKIphB8N5QUwGJxRGHo0/iCoYjsslbixkwIQWcJLIeJIyJ5EWt1Wp3
Vi3OEiKYGQmjrZvsJxB9zDJyogn8hhmMwSrx7B/0H3dBGX58gMLRkLUWL8OtVr4m
cUJpknqO1VWIsY0HfOvErHJc3q4JnSw7Bjl6UnrPfcGWznUHE0VSinUinEwC3nUG
RFy+7NISqJv6dNtGaNd7bnmVp45cqe0YDAvTxlyT2Y/0fGX7E6dEGHiThM8XNOb3
7KwQpB4nn1+DUaVoruD8gL33hTLKmLdQ+tnG8WhCQwvyf+osTB336gehMlN3mXBV
EguDiVKybgjRcZM1TjMNYqaxIB7FtZvkqu68yAhzRMqLlCbczaWd0+dKYlT8nw8H
JktIBJMuygNaBTMvqt67RBY6c4T78vBJm6TQjaGQcW19kHmQlU2hCiwO0m9gXuJ9
IRVZ8UFYj+/CSdC5TnRljE5ypKybmuQr0GJlTMQxxEA8Ace4PRVNVnCBgSPb2djp
8nCtYzQezRLfQmeHpR6Z56Te3nCw6BwWRw5rTWyW7aGuS2SjRw3UcZuJ7dR1bov1
lgwMQp+bKSkYL9WE8g51b4vnKRhqjzSUPUEOTTpha69tm8zJOHkbdZsvE3+IJLa0
Ax53eUiB/ZIKgCUImphKj+FeanmsdWyMEM2InUtmdGRMHJZmSlfHNS07QIDWCSKF
t9Re9Xxywo2akm7D+vopvfU5BOg8a+UazdBXMgc5fBc7F05h3rsqXRjgM043HuDM
vdvY664b2tnrV+zF802W5taswMl4I/BMKr4lifihjppZJTMlhYAoDssFwUePi5D+
IFQZuofhidLwxc7hw7vRsJComDKRbHIOH+T2b0lGjlhDnOL7EBDabZQ9I+Y50h9x
w2O32uxw9RHo2VJ/fUfTJodnI9ke6LJZDJ77YeELz0CImpFjWzFvx6qhNz6QjL61
ZlxfzTWp2CwMT1EjTx2mtZibJCM0SGrd8i/su1KcD+CrUh1r7c+k2EdYvCpZs3KZ
z02U9EvTcij+zQFqMp5eNS9mIIS1lnS0z7+OUYF1Dh0te+4snoWKSguyO7efMHm1
rvue43hUSzscJ0nSkfy6msML5ztJhaVHt/aBGvHMpPcZ5d9y1fZQAcP2O1XSlWpO
bGYw1MnkDbF94hTm8A0k+nIM0docjfhtBuWjFcH+8KPertrWv20nDKaal0I5310s
o8CtcnZMCVDr+TULnsQpM5RH/8gMGrXN+6dGiElbuhwwnn7v41w1anPwceSgmppX
mBw4S3X18p3Jybf1SPHgwg2++ZbdQC/oMWKlshjZga5zuBpdFVLHmQ04LMrWPsas
BbYWI1s9uw2x3nqMshVpeE/UnQU8Ef13pzcDtC2vJ7agHNd+Mkv17UuCy5rYpNmF
9vAFvqjYCDYsziFb8PbLiXatrur9MJqzujufG6q7yLMujr11hot0X7MexIDu5lei
l25yUmedRrUKFOdDi2QWi3RDQX5WOjd0ffL4HncPsafvfYVFkjkAExlXp4GtFONB
d+sbTBUVa9cnDFrXd4S8DAQVjNg2hYWDamSm3aSXG06DPfauraAlHJCxNwdvB/22
XMAAmah7B+KCzeO3J8YwyT2BeYLFHFfX5TYPsyQ72DvAr738qV5a7OpsC18zfng6
2TygN/d2XHs/NgyemxdNFPk/d1uf1fJZ53ygu8debf/ZTnnHoMjNPHgLB6zi0Xco
73Z/6VZ9pH35Jeyy4+OszqOXBiufJn2EcJPiY58hIlzaBl/AF4CyDIkLJq7i95Eb
p5guCvqAOpqQg4x4Kj0UwP0ecUk+ooePSKnmD0rnsVi7YbuBZY2Nw+sUaM4NL1OV
JLkAfmrdvVKCc7ErTRgy4iTRCvzmhFbFdpcr/mjoaiaqMWTVzoFJjXd3RtEYDZrU
jMBQVY4+tko1U0wwmUp8qIgBkSa+LXeIojFdCh6xhWZZCxywrunc8NhPN9u0EroE
QJIDc6Ah6mGtvtNgyFXxZMioCqPlPBvK+RGnbVlhdYki8LGYfERrxPZF0fT743I9
X4ni1XQHSZwp6UMwFUmQfU8kZDIPTSl5XTPWNIe7f2tmi/2sTKUeCGa3G0rAKnLn
Rksyw80P9M+kWuUNS37rv0jGSryue9MmfC7sozHMQdO9w1LvqsbM2o25kYcz4bSL
VI2fTCghdD6PKcxZey059TkYDDm+8pKfIqfmsONolpGq19mYz+jxpmjO3hrO9Eto
1nrCqMFxI5CpiiSlkiDwvn2dl2cVsiN/7RlwD0ZunjJ5bD8oifrdO6o8Qos+mJ7y
bwm3P2CyHhbdv6uGeWq2DRMYV+fKYLmCvwvPCs3HochyrtqkrgfjmwP6Cimc3HC9
1DDIWdyanQYRMsA8dRsOp/mJX9s6L51TBVMpAkw9hiD2pTmdVJtBwEjcC/V5aVGT
nTLcMf2Cfp4f3Q8VE7fyzwJs53d4+P4luUpZVlRVKDnFUDZhLfzGt0FPf3125ocT
qN8/9CwkNdGKZPwRNZktLnX0A6Fmg1uwhdGP/zvs8HHztuVbpFFEQawWJHHnkxx0
Qlq3JfQC/rqRs+DcWebjpb/AHIXkwlqokZBb18mITy97UZNSqTtDPFJLtx6oBGbW
0bIUH/8ODVi/7NNleMMsN6uen3TPCb+iUQorI+7XFuckMjFFMjl1bWg2Twz7FgDm
xiJ6QQpAKMIF3v6S8ZUvp6Jki0QRD8s+P3TVqX9rLUGq8VegM9B7N7rWmBh0LvXi
ocCsEBLJoeocp/sMM4JbUs90+V8BOSxDKcBgIGTTPyxkv0Gf6ClCcoQx0w3CDp36
vGqXhNE0vCOg2jfwx/7QPx1uOBV2/hoelhPvEuWb3KLDR0mBPfQu6CgHhRVmb5vS
UWXmeWgcgBNyACqYOd7kIfOz3riYAKZxc/oJNeAk8VTuVeVYUL7czqVy7Cv2q33j
0IfZ9pSSvKPeVqDFd/n2GuGNWFFwFoNk3hcA1U2N6RJlNry+QKP4Wp9fcLOJS3/c
0zEO7lWz3Uy7V+FDSQvp9xtd1EQvOh04RHa16lDAiqEinkMlZhihPeHwY7rhZgKP
9ggON+TQzC6C+hvkn4Md+ieki6Ecssao8wc9aJGq1m69HgU6rwd5A9FSUnCyPvIv
viMxkNvMV5CspLFbtMoukBOIQHvjzCPu2SGIf5DjGe+E/iodnpYfX4Pq4J6rgtFo
rg4Qbi78DG1SCqQYfwVMMQ1u+nCk98/WFN4PkX8t4sjoeJ+U79tDdwubG3RRZblD
CF2K+EtnvERS3lDuT2vNJWZughbW9u19ft3Ps0npor/p4ACdzfnfbibLBZiqZUj9
8i5ZbagWSN8wn7BZiacgfw7kLKKMuc9nv12xrV8nwB13jzE2oUTPD5CZVv05ELI2
NWJs7JaCLwAysfTDvMdiHKdVviABWjB87fU5WVY4U/20PMH3pXyiYXLC9v7EcTdq
HiYR5KUuVAUH9Qr2vOhdIenEKkj8do0qqfKi1s2WVcJcaQ29+qVjYm+EP54xi+2y
lWibLt5iqjvtebue/y7LM95Hj59+czNwr14BatL2JgqfW/fsluzjHu1Ry79C3cx4
4vR0QnTqGTksuoQYyOLmRnJs/EHH7c6DlotIB7MkQHFUxksmIgZ5151cnrN6BGmO
XbgpHHOubmBE1lJZ7f7Upzy4ngyZeXzjKmfOIrVKmO5QZenbDUp1D4MXjMQqpgar
w1uz4NTbhl4bz29tsq+UMTbI170FW5xdOs7VF+9tjksAUj7FxFtj0h6S/CE8ZW8n
kxWF9FG/d9qcFVr0uGVVjX1avdv7BXyUX5ZWlBAIDg5ZuFn15prvZOt2Rdd+d5y4
hYJ4pA0zT3cstwXHx2JWwRqjMoPZqSRhgG499jeAU3Q7pd2pfQx6Gunr6f0sJ6+D
MWARcZrRjq+ZPHt8E6gO5MUMXILTHGASFS4CI+muPDVPxjQbdzwyvwmu7iZuinCV
E3PuxTyrOGzKL2h2dVgdmUtOL0ErTtLnrAGR7b/hvQH2IfpczoU63MvXzM5+vkXe
1fEmI8XrcAicNNoErfpGQ8L4pJeKE52WFSx3IF8HeW5fiMY5yEzmSfRXa+Po66O0
ZkDYdl9iqERYIw2gabVOO9ds/2S3m/w0cRBfWsl4W3fKYDRtfLrdSxu5GfGgcs0h
fX0m81CApFwl/7mOd5nygbBQvXyMO0gz8XMmJ+8cjd1AtmZiDAxEMbJnitmwA0GQ
FvveM8bUtURL9igokn0p9lsaQNdZ0wWlAm78UGu3R+z3mjdHkHQaJ0OjvVCnp2oB
BtB4kfpEXG9oaDJEDLYZZ5zyUyQxibC1r64Rx40bsbryOmEa1TI5apoBjMgxChki
xmDIigOQlCnI1C5diFuGdL+B0KPAM1JMOkU2ocUSIZdvDistateDjxaUyoipB4Qv
dILlK/sVBb/X6r+RdtZCKTZqIb+WOxeinSvcpFyWYt/fumja9dry92c9Ji3GiDL+
KT0geT/hnN185tBCV09K45twDm4/zWq1vho+HGUgDZmruiKVwf0hD156HrUGfeco
ph2tlMnjly1otYXHdOKiFld2rCf4Yvyv/HDFjbl+zp7l0hVsih7SYx8VNFyQf0e2
cGl27Kj2EwRa9XTxED1BVWtXEZEBnfd3mwDFTpNfM1TVhHK2fZuR4qBk5uiMzed9
d6xz1KbMEcgXmAAUMIJFNsQUbYogdh8cXAfB9Rinpiamhb+tXFgYGR32PBZygP2d
uMbrvO25uIC9TTDlpQxEa/nGFmIlAqFhzGur7B+UMpocv2BLpEvi8Rc2R36nukbP
bqCye/u3Asco9VXMeWsn08VFwzeR0EKXhQfXjmWk2Vj1Dc9cPpKRqOSZq7ve0qQf
zN7MJzMVoVHEzKb8YoxEPdKR5lPKfCYMH38MGRbHhl+K2sVpaTM1qYOBXy9bR1kO
wHSW0KH0zCFUeKMXcKBfTORH8xfh5rXHL8z9lQV2hvRQWQWr3oIo8Gpg916R62qE
fRyZ4iHY+1WH429nL1KeGbeH1nfvP8NCjDYLyiqvqXQzntWOnlqs4uhSCoLjVdq1
WsKqFfvSmRjQdcVzIzhpdW457Ni/c0P086lqvLCG7+aUJ8REsbaqqzx352/uSzDQ
e55Tv8E5/zWRxS2x24CQJ9eFaXOnTrPFw4Z2kGqRw0F3Rd5zSQPilbRBt3y7BKam
HijEWaytFwAOoTRedWVB6TbUhSdvh3l7ZqtT7QyN+ic0h0sxrWSORP3QZlDP+XL5
PvebXnMPpWnPPKSvOkptwkMm3RTu/3I7YCWSf0dl6zK656m1z+EyRLS80Vs7hpON
feki6WqEy8TE9u22tQ5Hiw0kUPkPxbap8vLtrIYTOhisD5kLluOIxvmk1fqZKmWT
lsCuwDzYcDoUJjbOsZFm9+Pr67D8tSF72pHI/z2fWjjZVGA9KjEj8VWnT0zKn6GM
L3jsCOlIVO2d5PWI0XKv1+0cmPmrE2VLvIqePEqqSOvj9quieCx+Tg4I7nFTi27h
eDd69XpaA555CYN1jFktlEpk7RCZqFw6ku1AOBLgM84k8xj3iWQKjL3FnhPLgYxT
3jcRTbOeE7+uycZV2Y9LKs/gusS814h7JCAYvRKM7a/9n1QLXfMVMFKUM4gfZd8E
pjRIkPb9rn6KjHc4Zt4A/CY0On9uytcY8D45MGfMbME0aWU7o0Cf6MAozK+KHvXP
y4ibVh6uxWzNDrp6PEbN21weXcpBDucbuOmHe+qNCGnAXuwtMTp4AWGYhFASE8T3
BbwImL70cZUe9MBymXRmvKnxc0HmxDEtms1Cz4mJAHyRjaGLpuH4UsZvvnq8SUUC
06TvogB7zgF2uHHPl3UqTkzYchDVopmY5pnhpWijiWvhiIZIcXkr6SCo8eAV7za8
2PICxkx3AiPzU4BIhHrEkaROWuG1kvUaYG+JD3bNK8d0qGlDktRYuu7wC+rsRFMx
CmhwIXNXnQiAAnHhzYqVAFAz5MFV5i1lFqg3vfKMnYWTsAAm8nAmwW61zqG/aqhs
qXyMMSTtZqV25aATQNkbT7y2Lfnt7hxtOVRIdy2PMPGGVm3p+7ZQG1f4Niznymex
qORiWSVNjWQUpUy3Ar6Jo2dlzcJHdji+lprtVKKu87t/Quewjn5AJfli7b1FBi04
BHOz+6FvsAZt4/bMIEvyZmALKvqlKvWGKHGd2qw6pivkLkfYsRBfokvqN/tdfeuh
nkPEBFEmE33j9RktVvcqd1pENRhpO5U2kFxDoaLFExBAWe75pOPFUM6KjIaBDe7m
Z4En9U63GOFGhuO4kia/92GlM5aELVlKWX8dWj5m9ST58KKLwR0zG8QVt71/PT1c
YXSWmqIBJgkG0EUET36f+a2BJNkNeq7ivVo7Jnf2B6p8hReLn1JnvmPQh5d2AwKK
GGE+1ANw8P2/7jPMQ4meKFaVKc4s2Cw+1wVB7T74WDoXSoXNAZ80JvQYavG8Q/jH
uLtZlbFQU/f/bN2FELsRRY37/TIpXEivCIKlO3zYmUfhloreOpKpzC+02eoGuuHD
v4t0PFzMHpm/iQUSzKOEdafbJW8q+KCFWQwQDwOv/Cr+w6g/j6dvbhdJH+bYjdLy
N52MOTZngAe3Kja/CeYqkosXnGfoYHmYDg6mIw4x1YQPinKxnwV17KFjgwEy/39i
bwvFzUxw3H6EnzSQtkqKXnV93y1Yx1YNPeOU0FViewkpzwUnbbn+Cc2FdMHs+TSu
V4fGMttc73mNKNPEBvmdoI9t2Ey1f6C4S3uRwcw81iZr7xIUBL1zGMK8J7PUvZut
r6Trt99JTXCCdyWTmICTB0sMRKr4qLLYnj1BNpyxhTXVVHn3O4pDd4vwaMOfY5YU
1ShJ8OD+kmo4L7dliVoTnFTRQUTf4gbRVWmuOzm+aci8W8hYwzFAYMSqVOkaEtR0
u6yQXbaovnfXD0P0XeUSaDgz9iN9mPl70thP86nbCw5EWVxPotRuzQa1CEdCAsxy
J6eUReD6R8Afi1zYLSOug5NUjUP99ecCmAKNCgeNx1K1R6ncaGXFt6mEZL8nuoVR
7Xb+N4WQWsHefksFjcdMYx+rXFkDgd093mh4m22O5z49OxoMzXu6RquVXuax+aHV
7flUK7Wi2ywBQqdwZeUwBNfBfnWRl1UwNj5KbU3AO6dEHirfFboY/fuPmp3yQqgv
QJq7rL/lOaS85y6olz9zS1Pty/yLnzQJ0x1tUNKHuNPdsgbhxgD5n+Xo4Bjwj/2j
VAW2O8sPkc3SpYNxQa2gWs4qN/va66mzVTn+u0t0u585u8NzJmV0SXeB0j4Su2tV
aycLF5lhtOUebJ1tKG/nJuMtBgja5hofP+o2EuX4bOyMErsu+vVZEUQCTTeVX/XA
xQtKGp2dcWcMInLfaoVQdy4KgKW7E1cG9xodh+d0J2Jftp5f1doLxRcGE4HrDDeZ
hLFsihyk8ZZVN9Scg3IWspXoTJEIXbBDZzmyn/C1TOWw961TU0nxlSCpJ3FGaMwo
2XBiVMSXLBBG5PMMs30/cx5zndQidDrAYe82yt90WH3zw7ktAnjfDD3orfO2yhlX
iw1JAsVeui0He0PVZ8UWmy8bKf6ULJWR8DDJJdchM2sKgMcIWV/KjXIlodj5fl2S
EzdRcEK63yKYr/MhLhEwTaHVnE33xtVBqmN8EosUBCE3YjWL0ZvQYKe/isuOS/ef
mGGbk9VdZeFE1/RgiFqvlCgQ6b8mmGjgUtVvnPAoEXm6DkTKGmwjjfeivZjX3JPV
tWwg+BbDHu66WkMI2IzU8SwmqZOgGNWtAyTOk45hbt2YADyoisYs1tCaL3eE7wW0
OjA9lS5oSYyOQC+lnfpSt1+uUJMvqKbzK/uj7WAjikZIX8An8dW5UgVgyN/+H5Lg
MhQdKgj9zxGaZSD/VEZtLLJWlsL04KGSOogsRx34yYD9Mrs3fOROAUKM+//8n2EU
+YYt5MU1PpZIE/EFIMw+3M9hPvQYM0RVp4PpW2/QVY5TQMB16GkyC3xY07E7ZKMB
g4X1nJSj+t4xnx5J/4jYmvYLIR3fLKJPHgPq+T8wXixO41ZtlsBuyRLiPd9/jOE4
fLJU6VuMu2K/5gbC2kIqhv134d5C+hr7azIZiI2SFtazdQIMvkUfeFMkaky3FkpT
jhubfy8HXtQgqDVdxAHfcVAtFTs0F+r33CFzzdl+2oosbbUvqde06X0QN+r5Palv
bHh3D8vC2Ep1gTL4bwlZcjCH61HbtRIOtKqgZ1kSSVlAZ+8R/uWFDkGdUfbasyCf
rndj9dGXrM9qf6hR+8C4ZxDcTr0t6e5sjUxgNuZV3dBHvM7CZ13WHH6C7TBf9RrO
Y3Twki+wNNSNbv9HjlYSSkN3LLINiMWJt+API/jm+8OTUTgQEvHO1M682RNiCUqB
yooUc7Yc3dtAzQr9urnCZUpskiwYyudMg0zMcOFnPGaapePkVsaESgF7lT6by3sN
tBMv76zLPGsFjldWXaPBFeK+V0qAgA0QfNAuhvPQU7IbgtW1GHGavekRxk3h1CS9
4ArASe+kY947EqbLBJVLBmKZaoXZ8G6El2Ilv2ZgEha4Mo2rSQeR8HWeNunll1Dh
1SDt2OU22DHSFG3sm3Qw0OTm7T+e3XMFwQj0graO3A1fsQqUQvPI7KgOF+nabU+I
4uiDn3++MgnB660iRG6Co2KJ1BSHG+HQbiQWV6Y111Rx20pdqBofNosXBYSPdyLB
t6t2Ui9Zp/dXtnPBg0GXw3HqDhOVuxmZV9Yao6XQExWX2H51Cg870OlhrJIXCyq5
XWSYFqQsIVDS7R1FJUaQXB5gcco/+LooaNOarmkmbNZqhmsQUkZyIzn7cLhCuJXd
bCkqEsG14FNQy26Zmpdslvwg+gpvyFdUGQDAvWQ6nq/3j8Rgxds5hN4YYdVc23qi
VcV6xylgIqKP4gB5WMSMNCKkcpCmPVVuDDjpnhZBBtje7nXWDmcUz232dQawnqf1
+aLy3Byq8MJJHO4JxXD4K4M5svKk8fGMD/4nnA8lbVyjtgqhw/Mlbg08ehyU8s9U
lXOCjvYeBeSJ/OVPWCV9uu4cA9bbl5PB2RhwX6A61wP6hYSqd1zaMvDF84musl7O
026AE1jNQK8eIA+8Tn/EBmw1x8L/oJLHj2FGzqjxHACvWony8njDjUxg2lI5ErBr
91QouNhUE80rviFRN3Z8cU9VPBNYVrXmsLoioofIMJ+m8VEELiy72TXkvit1Qtzd
ywvnDVKlIzofu/Sr/qmRdCgdATQBCjjjl44t9dbLWiG1AI5a0bEx1anyizIX0z9h
ohQu02ZYlzm5d9FSejic3sx5vPXqxxZ9ESq2wBdQ2qdU8jYG+1P69xbh/PrueMsC
8XzBxtQMjXAntKEk68ueEHvJF1Ke68fqMcbtifdUTWDgf0sd6EMEKlHGe2Qpfkmg
g9azgAndHL0fHPqXamr0QeP9eK+CrOwtN18UkOM12+VGn8YywFYZ97tRQ1GITiAQ
S4eUbBFC4N7HKH+Aro0SlFkZlFTFldcBfYoMzzNTv144HV31ZIrzpX0IJNh1TgEn
a7NVipPag/AS4hQW5Db6/j6wgvJjsaUBcUGiI3BnZ+XIDFFA2avqggCwxcpPNVXD
tnD7c7Jrc9mEozCiQCnkvMp1hC5PJm9Ea8gqtFWneUaJywffkzYplP3E14YxL6xE
CCV1GuVoCvIy5FiQ2a08a2Fo0f0Sk5oVvSzbKUAU+wyI5xGF0TB0atS+YUxsdZB0
2LAqXtNsBSlPWkjrkcFEJYWgnMbrwUdYTE/r3KunDC98yEPUXTbsZTtINAFtOvgo
/v0Eu4ssh1Q/mlUvp+Vqm7cdP1CZmjiEci7ZVa7E+g8RS9thiD1L8qmdIposYhWj
qDfy51tDKzJ2/tNdv1rjivKt9eSxbKQrnAB2ow4lOp52ZTGaWpg3EWOsEgpJxopN
a1PR0oTVuLDGOKlJTQvP+cpdw2Zd3LsXijt01Zejx0HbapoRqglPDYsDeU1tA9xC
ZUMnFJ2X62JbZevlOS/jUxYt/EASAbiY599o/nI5N5vooSAcoxAJmGHMe4nNmCOv
XEVlasj62fyRXx8YGvB5eFp4JQNX9xvM9jPdZpXVXSzoXb6rEHHaV2f+GKUFNrFt
ks4L8P+L+DYIITng+NtYYZ1bn45DaGp2y8MxSyCGygwczO1AVHUjp3X4IuqHHEZB
/B+VJs2L7D/2SDKryls1J7qX4SxB0oc+rVwLVc9fyqJgoEAd3KP/FNj0bM0oUEd0
gLXu3qRly1CNCPAW9F5Cr7Fb1xuRJM5Nc/vSMPhPeAE+0YzfzRcXkTvjaG1N2CxB
dbHEUlVQ1L+XJ/d8pWgEBamAcOXJGZHXVHnrl0bTENHyH0eTAxaxgppRXTJ0ayC8
r8ljvXiWgnBG4n1ATvul5pPbg/UUmeBM9+WWNIb+6T4ctbhoqzFF3+DeHVOTT0/y
Yopi0YtsLArj+sDD2AacNS7612U/rBG4UeZ4Ajt7+6+IO8qylF70+gh4VOflo9jN
ae9tNBI3GxctfrvZomDkCKTFJuHj6GplP5ZFJw6OENf1qLpmW9K5L5n2f+Ogdd+W
3p5W78oYioDf8EHpe69gKiVX9D4eQveE3w0BunWXzT/QK5ixW9g+uQVP7HBTEpyJ
pM/sipRaKOJLExbZLKNV1lXxKp0pyXUCyd3hA4KwKWarc8+Ols4xWjJHSnMrjZ3E
cDdIzEmyCyqgd58TqAGJk9/dpgu1gLuIGquI0hCdulW+I0af0WJE5i3JG8TYdWtS
KI7i5eSkgMEmMeRzZZJEaQR8vjbj7geOKsIe3fmgQ5mMFQiesSPt5lBJv9uH6KWx
W3UFYKNOtHfN7Ley/i70q0J7Nvl7QXGHqgJPyDfaFaSo4waRhEttpPGn6QcWlA3t
KCvYe3fltsxWKIzExTEfiMCPe/Af6PGLaF/OrELRzxkxAtZI1ez2SGuePNoMwxj/
gzJL0IsXGmae9YUq2+/WICfCbluEJo2MvoQ3R8ujWptGSpPGEneMSi80L09OQT4L
JLIaT+Ez1A+DbVwzzaB66eOJ7nEZmaCWUMpGdXhXFyhQxqeVVME1RTh1RLY/h66k
mYcO80q1V9c6cOnHAuhoZotpJmYqwqHhtJEahowsEko+Y64FIz7LOPvT+7mhBg85
BeiKrebOGwXak6ukJ1Gp8qwFkuJOH1wL+LnM3NsiuVXCQuqAtR3I7ko81jmA1zZf
7kBiVlF1t0HAdZ9++wARvbbcJaYlcqBhYSvHJLffyssuywl3DuX+OxrCun/z7E7g
gbCnTMHm+p4J/Lde1jm8z9dpwcs2AGqexpuaYJZyQBS0Q54CkOm7S0aJNw1OxfRD
/qu7kolPxHzi/r8zHVh2LJ/FTqKafHsN30pOJrM6Cmg/OQsQHaEiISqauMDvBITp
v7GQzACw3qQt8SddFpCuOG3vJZFKxglhXQEs1IEMuJZHOJvugdGHhL5m8Heo38rf
armrrQghtnw8VGFLTcJ2KiL90I+ilca9vJtdPGoqeHb0/bPlWbBp++JySiQmLv+d
Qqizlqdrac7nbhXmOlYMccZpyEUxqoYI1lzisI+0RyM=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NoW9rNLozfNG0ASTH4KW+4SZv0xFwwO4yzuoTClwTGqTYu34IIbbUjlYRB/0+aWo
V4CWpECYaRD6XnCfT+rWmiWfoeGC56LoA3wYrRuQFJNRvrVpNq9rPydeqNCT2yWu
NL1v7FxnHl2Kq+YQKWHdS2ioj6fKEa6G/iI3/i1l5ZDWTP3IiK6WfGYbAZWgf41Q
365YYa4Bz6wKV3JiHw/xWeIUXA3Q4SeG/mCPNzJ0hV35R78/hRfTr7MjLGvxz0EW
L3fEKz1LT63Rn8nxUZjVcvlw7KY7WbPlgsNgUG9fn+GP3Osuroe7JYOyNil0XtjH
hpjDi0GzoihzejoEyQd6Hw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 544 )
`pragma protect data_block
uNLG0hUWKaxlyIdRGDx21X1mkZyrzCuWeoqXjb7YpKMqb/iytpGJuC8nRunYL1ez
11GRn2JbjW8W/8O7SPGPM+1jAmmpuqDNG5Xsp+4kIiuJoE6VOLphkbFDM07NFkh6
/yLPUdfNi0x3fmyt9rMTfDIW1X3/6rqDlu6Sivbx9NC4z4jJ6z/sU6e95/tUFy3Y
1OpkQQX9iDP5jIOu2BOFxEx4cuEPFRh6PLcvp+6vuU0dP9Vkn6l7tjL91vNUCti4
snM0ZEgRs3dzDHPWHlzaPu1Y6T01l60o+bI7GJrJuAPoT17qVketc1CdoDeK940B
c5MclXgQpZ1gkflRlwd6RbeBLm+H+n54Pnc8PiZ6D8yYnrdmhG2gt7pCG5JFoZeL
Gw8H1NjytRKpeC5wVNDH02hevYurNMXPgyQVggmJEwR2fE40ImUk/wUssiM3PiBg
nzY/0fjAOA6LVkylkDDkT9XUFhMblv9q0S8hrdynkjxL3tBfgd+EivUg+jGOtULo
mnuPhud7FYzyUwWGcIfg3S/YTMRIC4AsCue20JF2eSk8fKJGZqOMsg+gcxOVXf3L
uHFXcNY7Q2Eq1AqBDpkMcj0UOl9ILzyTA7yRACnDFFZZ7QUhMexKMcP8HVWEQGo8
PIUNUz2oYAW7qF1m6rSWt/Kg8tUF+IgYC7FWyFUnYhx089t1moH8iDbjlYdsBNcP
iv7/FqAcgyriM0Yjuyz3ew==
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NTs0wl6NaTYtw6DMnH62LIubC83BFHLnff1O8mY+fKYC1x3fZbaPxkJdG82MHeqq
bPGH5tzociGy6ebnqIlNtCFAY9QX7sllz9Ta76kZSLwStpXKCXoxp/EE+rGR08W2
JrT9U5PlbaGNE6V3qLDLSjB0o04WN2XPJQOzw2o515gYzELmKlS7a21l0EBJMnvK
uU3CkwgURuLEnd5ulqrH2Ka6zJ2kyxmQ1j6cbhsWmT7faXbb8f6D1mlMbB8hwVyo
BiqrdHULKqX8jjGflLEgEy2JTewp/AU3azEWX8l9x9eLUgk6r0dozhMDsr/D03TW
IRuiF7JXfojJCAAuTSzpmg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
0LrwzEY+YQL8xU2gZSwAXX5YcsYzI7wpoDV3zXVZk/x3b6j7gFb5pz17rxwyNIsY
tkDhrDuAad8mvAmQljeWZGJWnccvTN/zDGX1qk5BHMFex9rS/lBEuWHtOaPlotv3
CMQj92gwMC4Uk/s35XCfIxZL69eh7cqtR2WJq+mtBf1XLJZgi1cbt+tVbsP1FPMe
JoEmbE/6xYYP4gcrajgyiehl1s/fIpisAwFNHcQr0lkApShA3JQr16rzjnXd/MT7
kXhbAtpOAmlg/niujyazRSy2H70kqqAm+ZXl6Jd/bn0u4K5n3batcQoqoLk8i3LF
DD/XbXZ+63XB8/WFwSCer/qlBOjpEgpC+hDchnziJL3OhjAXL4Mccmu/J8q4aZzF
ZFCYVPg4v572qIpoDpByy6nQRwySuSCYVGJnCviyBDM+7AA/X4qAXSrkWsbmZMU/
T/FVynIGY2Eve725wu+S3slLbDDmAelRa9fEz8eEThJHhdQ6ZrxpSDgFKRGsbnvw
NXi2cqV3DKlSkJfoQL2WKJgToqYLTLxhCNhK5xH4hR9wlrg7RNgqngcR4ZIt+M2p
YmZs5vIUj0oTKz5wlqzqA9rvTwlLW0HLcpp7TgPn3Gt2BJUI2eSPBgYEMctpu8d5
r2vl7jncJ1ItmOpI4pMMmdmrGmDpG6Gfh4i0+UhzMrI0VuFIeShgTEOP/gxDlctn
7UrfkZunLEFqaDS04Grnxe68WJO38SZ9yOF+hjPIiet6eMcbxsRdMJV7ang9W3tB
oqPwBDjng/gcLgulXaGDe2mPcAXP5Da7PmlYJk+vMce5POV94Znar4w9UuHGP07y
lypyx++CxqCgKI3bdWSG6p7P2l0AxONgI+gSfUJhya7ZIPJGZ/mnBT+7EAf7zTO6
6xUmqjcUrhXK+9s5au8M+D72CsGnv/yzBm2EUZ/HNeQ=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jylntsAQVqai/jJaGL3KknVkTYciB/UOaFiswlZArtVF5jXsfEYrxdNlQKF2C+ei
1sW0zHenIyYwKRWS47jMR0+fTimTDrgHetCl5XR2E7RVp/wcjsRkJJF/jjiBXHr6
BJhVF8KlGybZ7qoy8bq1WkBNJhze92tcsHS+Wbdn4NfbgZwV+xVxJ+RqjNugSCfa
rPgSqO3tc1lugSL2zAkb4gXQtyPvYSMMnL2+wuRzJvv8aAbdUg+i/VXlaD2MnoNQ
UYrF0gG3Ew4lwnXth8cWc98xgoQh9EtJIRqYF/6FBRkPdW2lmrBoDV3OsJ+EUCGb
3bf6mVcdzlOUutx9EeYgiQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
KddmpSs55Oo+odiYslyfopCtVoAlgnMfrjmYwTauGqsUZLBgbutSgiVxH55ae5BN
/CAger81cbj4nRYVNhbdpJvGDQIKIpEqT1nVEFWlXqSKSOfZF+5Lpig34u1cznoZ
eyyqZJ2SGmk2afIq1DqV7L6MFEHrlv4JknxdoWBJftzZt5DHZnpLawVph1BzKOxv
PFkcYB6JHjvlaMQJvepyuiqwy8g7RTiXiNEQG6Io7D+lWMWdqezuUErnnjVc8VTP
dcUmJp1thxfHalK2IwrKbhT1V11plDqEOO5wj6zbCFbY8Mhtojdb3m5/tB8fSXYe
QGsGbMe4rtsJa/9Bp4v0PkRvsN3uLPhwgwCb581MzqPOBaIiDHUUPEq2IcWKNWqr
BUWO2IWVq2TfwSo05TIklGOmNtKyL0pUs95ja9WllYRRj2u9OzOivHOgG7MhSs5X
wahX2CdguCubsHlBLWSggrwNal/Wd5pGHzyGpVWEUlVVi+miOAAZJ4bKMV1F4tun
LMce6JOkzOiiGj2Xrue4pOqaYivBjU2rJ+6/lwvMUNKnZ9DNUJNlZI2ho+JcBYLt
TUNLIargWEbvqJ207QXG/QMaAuEcP5YN/Wcbq1RLwdaRVrJu+YVZ9otXebhMErRk
4rARYszwC069uch71J6TG+YRdtY0hBSpZ+RBObthCrN/5lBuXxMUn6y9TSUlfqJk
/nhyR3CXSXiCVpCSVlRj7Hvqs2SM1PSgilhgEMyOpIZyMkrkIeLM/3uzPgw+zErW
0ssp2HkWQw6LkVLVpp+d58MXGbj0/EoQwWlJwv88kJ6Kt00SqmKuYPUj7Nxkf9Z1
lTf/CUuAUiSHFmfMHIMomO80z1QGXa+wcm1gYeytuFfPXArqd4yzDiFMHAoG/5lB
ko4RvefkpctPGJ3Sl6k5HuEEpwyP/6hTGY+kQTvfcasbme2lubivfh4cfcEjtAAz
f2kNvD18Yu692AMGzsut4yWZyA4/pCyDZJb5ibyyVyt3fpE2rOtFaBXcwlBnCjiD
O0d5qkSPhGmG23a1Fs4rMFfPo779XWDR5QJlY4VjU2VpM9/4gt8A/DmZrAG+v/9V
Fx3Z/iT31CCFSnP9HsKtk5vvEM/jL3QXxPft4Tm8vLTiNYaOPoKl6K7xfOSeB2D5
hfXMqdjYGirEbt+GoOOFrM8JMbvES7lMshYSd/woEmTU5qaP4Hfxvc7dGycxf6Xx
A+IAyfy0LjngYyy9YnNFjb5Dtr2j9nrmBhwT7NQO+Q/jjLREWz66GwW+/7oD2jkw
NROq35sTseD5q1ev1BwiJIjcaeG90rWIk89OTGQxNWWime3RkAqnwb9x3VIQzwtb
Tx5J+V3kWMvfXeSWJGkx7F8NT/MdE/r29jZA+CwcrG/YZ8gWuQQKqgrQ/ZWHByUa
Z3aYs0bsrlwBeaUZkvFeKTcCBIBHdFMHTaYq2ctxClNfZfN7KTAtmnqXVOhff8XO
G4ILFcIhSMU6X2pGmVSsESbEUdRGqVuiySkVqspMoJI0XiUrwH2OY6JPwOzkoF0O
gWW0E2M/TyYNMAPQO5kMsFXBRFU1g82NbOGqOhP+d8fbNFIP/8QOnMydQ82YgDHv
dXqYKE30T9yrGWYmtI9coE6aNof6PykucAlLTo8BfXv1gRENohdXjFKHla1aQIEj
eDU+gf0rDqMIjme6NCO5JbBdZoYwEN26gBAXQxGX1sR2RtNV4n823VKKmNwCMVvw
ipqws3SMkbc2qO/EVnfDztXXnuQDitEYoPe1wnDYbj1Ck2XpjiaCL4rtxHKIBVLt
momEgVnA0PQDsAXS2ib4pSRDwlZKpkWm5SadsTIU2mU2rKar0t/1eDdSSc2haQr1
Pek6qJyiwl5+oLVZCWMSfykr5dHMcG6icCVvtandG75zSY3m+zUMCj/9//AJKbo1
k8m0i9/pdoZdbuQyAPwnCWljNUZP7YdmbkSgLTjqPQTYYFYICY0dHPJ9164J7Wbp
eMgjsBsuh2oCACklC924I2U9xlGXSpNRFZOyZ+C8YRqlSGEnSmpSJUEjfufs0S6R
WhnDOLNjIsBD21nNUVOhpBG4bKP0V+F67kB3pdVe/OVsb+nsmDuUcjoxlGI6yyIg
WUeuezidD65QlTKz3abTXTDGS/7ww9N0/2bi6hXhksMrSw/HjsxJTIZVZqW5dJqP
hDLhU8TEHPYhH+pfJgAJaOWPM6DeTuTdvuWdPmI0BUeRh2ZD6btnerHdxYsduszc
czR4fH1xefwjz5ntMwYWlf8Q5Sz5Rtqp2i9w8CdFOFSzJs13W+9Pyzifb0OK4wmW
yoZNjYBRbLkjLchL9ThSstoJTsSmqQFzEPJPM6WMpmg1oRcJCQQstSYKUJIh8C0Y
6YfsOOvOCcIX8kzPPuys2mlWhaYmDAa8LVXsZ/PZiPWU5lTRv348F/HWox/+E8Fq
saXUizewkU8pEc55q9SXIyo8c7K/PbD3sas/6uHETx+2UI3ara/4rWnquw5wzEia
jUP+2IagWaQBlythn+J3fyjvvr4hb490/lxQGAAGFsl86VLnFS8ag9W7k4d+CWvD
XuKvnzkWY7p4Jii1wlH8fQCvZTi/VwZNjpOSVkEKsxJwsNUyV9zAgr8W0arY5F5q
wd4/4q8X0J2fN4YckisdAO/uT3j1crdfXCNhx0iF0abmyn4xAZWtKmiOxWupM6Kc
KoZ/uQ0redOQ8bfOABu7z1Pqk+ClY8ipGIWrD6eFMdKQdQ6n8qfP7yguW2nNzpQn
RHht4fIDB4rZnIdCLwbsVHcu+YtItlsEVQeOlhpX2xpm7Si9EafePYOgb+ZdOtlY
1ia8MJxHMEjb8jRX5wQ8fCsFdXZJ7zGzlN9Zdjl2TkpZHCxtY8nkR9YHITztNhA/
E6IoLrlp1xkE4TZ51Z+/rZMuyisjrXEoACCauye/TmqoaZBgobkEt92Zl0K1ODj0
aN9F6TA9bZyOfW0EVT3xTi9p4Qlu5bbM9Z0M03jGJjzmp4PGqiJ3UEgIzzWBZeEN
VBPVC6gObMKWEkHOcazrY5nZhYuKPQgnX1gQJVHAp803aQlGUGJ2EtysX6p8/Q01
8tw6vRuG4By7ObkQaamVxsqBeUW+uAV+2zfwLuT0g2v3Hfe9aLziqJOpKqaRz7TX
r1gWt/jRGtFkgs77RcbxIv8JXlt+TQ1S94gjw9wiMboCqHulWXsrIO/l9GHJWSpr
trVpbcQ4tztBFt29QxEpDilEa6W45E3saCOhg48LIrSs8e4oQgK/J8vBhpBCQybj
7QXZ16cT2s/WHLwEo+DU0X3xEPMYq0LuKGH7bA6DDWryzNSVwh/29F5Kd+HCcnjw
n+Bc+RTFW4nFsA2XM8AwkR8s5H3GkRWE3ikcVjbRUTmyn37LrBT7B6IG75RAdI7F
HFXCPCQzrWFqTA8WipmVC2cvrVyJNjz2MM4f/8jj1WpyUwiVHqAotumAEVrCU9D7
rDwUyXMpmBmZkFs3BWBfw4TlsbdvF4afn7vKKmFZCLMpeIQx4hob3QRa7uaTROqO
zjweAiQVuB1s0dWx7HqroECoxnIdTsme7tr82Xd2c/Tro/sjI0tx11edqQe/ZEm9
Dz2/M15bLPvSQIj2NCs5IGqdqjvBV3YYXf7RQtBWrAckpldaLlLq5j3E72sT4P31
JQpfWyJlV/kT3p0Ins5gOmS7of7qW+902z5lgr1PNsqBw6dlDu7uhVyEn20Tkmrq
rF0sdA65dmCGxB+Jdx9CWMw3sC9QUHGOqSg/RVIXe/dbvbOc0tPzF9wU/jID6Goc
CcoIgxhwMfCA9xTRnv+jl/KLbVdF0lXdeaSvavNL+yV+Sxb1HeBxf3wU6xY2DjcA
FyoUA6lgH/su5WASmroaCpq+y42fosfrOwt7AbhJJd6RxWxTY/Og+dmyFiMhaaLH
3uE5QMPd5vnKE/9faDjmMbEXX8pFkVh5T+5YzQzFwbG7ItLFOIHdrVU6DITMihYM
F5fWYFmRLGcvHtjjD1v9Bt/tQAtn+YfzZ7itgU3D77E6lFGRl2G6tuT+PNMnan+p
gckjr03LH/HV6eB+E0u8lxGBiH3lKAV7knu0w+nlHsyfjzaB9f1vGeQWjudwfNt5
olRRqelymG4TMF2VEiVDan6v1cEuhj43S1iZAGqtudruaNYfLVcngKx1IxktxS9z
0UG96fPsqUHf0Q4TeVjFrHvippysYdAXJmC6XFHfkRdIWDGqIQCtAP//MvoQK2yn
u1nYvhMccTYOcFvit9+Lr8nrGBT3KkOGw94SvdD1yJT3Ne6TKfgowXQDoPMDs7Oq
Y61UoqG1s+xyqPNNPJ6SxesJ9TIPFF6F9Zx1dt/hlTp+iF02rO6rzm+2ExKZ6xbN
nQloXo8g/RRMs1HrV+897YESz73A71OlzGZTIgT3l6qpRKOKSus0w4ZIhi3Oi+0k
4k9oFFjkSBTrqub7DafU/38GYam1LlIRbakZD2ka9tInAVMNwN0hmNIV5iIOYgM3
0EMgnGB4QKuaoS+j71ZWDP1Di6Uz/L0x8P4ldn/6m0ApsotDfQ77zLxG+OAimdUs
dNrThzpkT8Di79D/vzr+EnAPIN7JosItisoTkC9yepWIhj509OpeiqTnArvj+85k
gGwNHcW2LbVzuPZhoCdqs67DRt7ckXxluOerpUsHutyW27iVxH4WV4Hn/UbwnrYw
fAKSjzriTlGUenyZlKLmmroYhWB4DlV10a0hvdWhnpUC2LFfFRdVub0I/e897W30
PRIKV+O7fjD37WPYlbj8OJkthpo7B2ypR1TPRidUod0AcoJTd4zWklNT0OQfKB9m
6z4pGXqBIfvK2S2Ady3IG+iAbFwijVCqNt4vFQZWJveIAcW5hKMZ8f5a1W+s9m0r
GuJFgoUgAz0cRj1DA/7Rc2ElZWfA1HNmPlu6ooJ98t1E3ylZKmXbFpDKtqpLjB+I
REB1sbs3P7o2FvlImiWRT+6CIHg5fYTugBTWDIrSW2JgtK2qCgvxLKlaiep1yAem
beL9i68RYXwpSvX+l5/eaA3QC2E/DaFkqw3ael08TiegaMPbfQRW87Fd/ci8E2/N
XfeP4noSeR5AlzMeFnzTVKuW3cdRcwSx8LpT4g2ZzB0SEp6UvkHF0ARjKpOBT77D
4HCOvEOay123xNZYmObrNYewJbsZ4ZsyT6gT5bQp51jFTFv7fs90PLHBRvVr26l6
31ivGuSPqeBMGfl5ZoUfco9vTiHO0f3bzoxr7b6IIubNHFYkOiaw7fsFCwjgAJFC
2bvSmYYEx9Qylk8S1qmgT+23gHLYtIl/KYDT83ETtr+eoIQ88834s8dsYugSEPz8
HBu4kXObBrTMGbdvDJPPk+b1DvTDj0svzDVyuesZkgW1jjAbUr1zksQGsOsSrRJz
5PUvAkjclTr9Q1aR8dZs6VJrv4UOQCm9st+DWNB7BUYt/Yv1WCX4yQfa6GpGwmK6
hL8eUBxXLN/zeKf1zW+MkHqVvE+hnveljOSggLO1tJ5DBOgVuZWHvN9ah5eLPdpY
U65taxSD9XuIibCqO6SNFsAlbtg4o6/iVzoNkB7j1qXp3uoWrPkUy4c88lrqqha6
EHdSSpm5T5qLfOFkC7fZmk5deVWQjTAcfmYqhMuBf6eNuAMzG/PGlTCN5d4bZGZ9
lRbQ38qzcawCeXfVWjHuc8SFal0z6oPXofN+tDSD9g7RbptdlIsoYFd9vf4dhaLU
xP5GTlYkPmw77fYdqv5kA0SKtKX3IC2/jEAXVgXF1NuWJ2uA9K2E6eEqIykeheUp
+tz0J3wqWx7qmWrYus1rbkW3nq/1/cHx1+grgw0yJ/oVlMUNmS1sr4CQEzcKn610
i361uMT3B/K5WHIkqJRjBkFPe1VwKmINiZVRMZHi504zgHmq/W279/2N7hnSZPgA
kewiD6xRaW5n46fGWW0B0DGrHoG8vs0vohjv7ts4cgTpECB36WGDtWgG/epx3KqQ
U0Rv7c4zffckPJkXgnYybjo1wlHz/vCMJr1cmsm3gaIdSLuQv7D9adMbO/wdu4wt
4g/mZEpYMkx3BaiYty6nM61Za7ghBMpJguNo02XV8YySBevELRabUzH13CXmtzlA
3iyWjgZ6K8u0Ca9yHSin4MgD2fURuRLZGnRLs9DzZIPyhCy6Mgka7rprkxg09SF0
hRXDbhYydvwuHrnBPDYojnBBCxc2/URdia7vfwabn6Jnq1aLVqBXvckWuz+vIHL4
xD/5A/UDmN2sNSk/urtw6dKPNmmExb2+MYqPJ9P5MXzVOspDPfmvVHB9aq5f5lTC
WQjMLtLON6AGc+vFiNxLBqM2Ixq/Grzfkl90M1FShJo7uv4qy/zGCF3zZ+0hBUBC
ayjrkToh4+yp/cqth2BFiKHRGmMPJq0vGbf/rM3pJRjyE+6y+W7cghcQg5qR6OJY
hDOSDKBQIwk0xcduzl4GjLQ2x6lDjVkJ7uuunNP8u07ZETUZ2+uQfmxAM5t+A5RU
Wj6CebaOh2NnO7WqiohJbgRwmlloddu2ag7g0Thh+0KS45fjxliKlCSazkqRfDAw
oWZuBE5tZovMQRWBkauo63VHKE2eHZRaXUvErcKx2mWH4Qnqqghg05m7iTrzL/al
5yNr7D4f6tQ7nxlayphc2qbj/9q8Ep+r7eVRcw5hCvICPX49i27dHrMGBI+nadxU
BlG1+1CFVvtxlr8K0IMX7TnkrdrrnSR+l3XlgzqU86Xs2uFcgLkhrUEMFMKI+SgS
am24P1T9eFw+0GO32283pDM1FTvvaQJ8/v1j5jyF4kYpgZegCdoWCGZeRTAbgbCm
5965Lrh5Q2aYz2VQvE/7IDAmeTp0STtRiJ6ZfBuTYRuf5SOfHB1oSYQVhpWh2eoz
G764Xlb7i0mmzlmhBYUBR5ic/bHQAq8GkPKBhibecx9rRHxglCUvDnq3I61ZRjsC
3PhwhY5oF9wjcoRPFUuIWDB5/TGW2UzrcQQsQBmwOTTnGHhMFgx2c/YTbkR9J/9r
1X1msKSIbuxxdmEggP99ql5GgmaarL+8iZn8YL7yDG6qhOf3f4jT0ByoiVY+b8Qe
KPCQKNzWLFxZifOJwyMns118Ixu5ITZpEJ9Kd4m6miCYnQosIaspd+w40ZEncG09
gRjje/JAGppyybhx6YyF31GW/ZmBV3qxIM7/47GH/mmNCIBE0s4+Cc7Mh4+WP7De
3yPmYuIPGZAp4YoeCImVtm/sdfTGIbQwZclU9KIqOZewAWtw9FvA1oEPAyQmKq+/
cXnpnhbG3f3aawm/A2EgDCDKZO3cb7isgHSXk0DnddmBDXUKai3tzUUN+ENTpQCG
MNDEgzf1MrPqflddpEugpH1DfeCBpP6L/cy6zp/xuWqOjrAwL3g4fUktEvOXrsbE
/K7Lqz/iotpNLNTQRnDClIY+/UMjLMG6BEuKk+Ytdt+MzacNUV8MvwfLEHtdMmxa
niOBPA1nAmhgJ4cU8A8Vp1xHG3ENLkU0Rer/48qmiUKxmviJAw/DO6l61JuSJt80
0GL2+I/3KlJn9mwamRnxjz73M2o3B0FlNfmaOQ4G51YNoaSfUrVzJUUkdkNUN3Ii
GraE8jhyNxMI4J7DBpg8Z4e48AVjEzdLrmWKWYrcTh7sqaB9G7SQNPg2jifFOXLZ
zk5IhpmlSwQ9oOgZt6aHDEihCxSZngyCtDbX2+AR5XTt+iGec9J03a+WOKvquwpz
gE73xyIjeGTsfNGCEFjG/TZ26oAxeFbtT5mZd4ztz1DoXAV5htV5w0ZvD+1ZlPPd
tHACie5swsbR2zuXMIm3JEWs8k2YYCR5Rz5AvbJOJFZAYbQBUhWdR2AkjIejd5Pu
g8E1b4pAqkMmijgrN09JZYkFOn0v9+xgcX7xdKdnFukJglm3+BnMfKUHE7wkV49y
/KEb6XZuPAg7QiW0Bmj7eF1M8h4YezwhGy0cV8sY8Y2UR6Aia8y3nBsCbXmXbM6Z
judlDC4dus/IV6S1UmwRz1mHMA6vu60D0LxESQk2Jy7nnYphYIpdXWN/pU1A95oo
3ZFcU6qW9SL/eGQF14sQTZ/2Ot8eh0+j9/A3wmZ5GkVv7hk3Qf+G18h5ev+eAvH2
EuOYIaaDXXqRj/9u533NulRQEjx3NUIt0y8vw3EzlD3uWuClv5WOHu6U59Q3MuOG
aWQ6z6zsQ3x23BeDlm5IQ57iaVR1DdwNbu4xEj8tDRpurTLKtMyc+fGhuO1BPkY/
fTx5uSPypqBMosNIwF38W6+uJW7dC8Kdcjk1EsnaX1oO4jQjLyt71iqYjl2kcG1Y
LDjKrVQFR9OpC7l6NR1lmm3lf4jX8aFKkz+HJ4l2HBXX9ng5zUvGdIVAhC5XE9YL
Z7ulZcZpYzBz3cXV7eMikXOSYiDQxf2YjHe1VcYodclL/Uo3WKzuPdrMIDo42RRt
07I9A0xh+gciaQuWA2hTckkKH9DWjc/dRFyCVP45iDAzW7m0fA5QuLTWS66B3+Pt
PmMBoRxdWBWLi9+kdm0UGGmO3zqJ2J5J6mjNErhsNVrM95yeFFNdjHzGtL3T9IeX
vEbmGg7WLYWpd6MmTQujUVoid5gO7TrR9NFD+QpaBVG7aDKgcdGLd78SrGiNFLRx
jww1/dlHSa2dThWBGRQ9JajzzrOWwchR7Yrxo4/Cod+EaFkx7c1Cz8YUWBERBh3F
gMbMdvGKWY+aaHzM1OsNficoslxwM736Ofk6+JAC5KURu4Iv0u3ZVlY1xcUPc9Vl
bwD4BxhkhXrRLcvHoA56ntQ2EjeT7bi0IF9+4GkPCbRR7/uXCzEd6jw4RDXkRprU
Y0nwkL9Sb87nI67iNpjViuP4yqIsBeHeF6DiW8R50J5rMIXEHGlMDPxX7QQiTNOy
xpZMAWFWo0vAdQaN3gM1b9+bX2gnQBAKzcVNyMUWsKPQMcR8na4HqrnhUbP3kar+
KZozfosyRDeijpVDep/3mIhVVkCqru+zbx0JSXu5kqDKQ5705kt7SNYD88B5NU4Y
TatcHSM01zXP5O+Y3V0tvFM9yLPr5Cbv2hZTagMAwn0/Xhv28zHYtlsq+lQ0HKI5
9VYgilSfTu5sG4/82uDCaygdHqPrstRPxcmkq+J2XotykYLiZ+BXdyZxkPEYkqHA
0QMATkFI+fwwEJMTvgq1OzCi+bjnzEqVMnmdRJshdaGku3qZVi1oMYHRX2Ib051z
EVVwlHB+h+/CyEB3wHZG2c7NLnmEYIqREqJCNyiaUaWisAoPNjkHyirlsE1SpWig
+eDmzGLl9XMVzkCrDDLJ9rf0wOawykDpnC0H4bL44tDEKo/L2gYw4keas/bzryzE
ZdRcM0vLD71+k0FPXfKFycAqzVum+B3/YhOjDffIhy5jPY5J7l718/cDfHv37jg4
8mQaSJrt+xIsHtwJCmu0gew7oEWigtcUBfpHjk4KiO7lfA8Ru2O96yck5eOth0bk
6to6H6GAlB7Iv4FcevxKforbVd8J1UVc7sxuzdrXboaHRz2T5x/pgF4RAPvViPIw
Gk6KmLqTEl21wTvFvdiek4akcgEXmB0jYiBzyInJu1eV51NEmByAgpPbfwouzlFf
36DymiNUIa7wITXHhMY9uq4RYVWBwn7lJwnux0NWXesPN5wVlvq7Qn/kyHrd1Y3m
k6osbSWRBN4AbEDNNjBvZSkTEjuGiWBX6kOvf9gYy+j59IlBEEC3+Xwxqpd5WjfL
o7LCcopK+tbvgoC1oTqT7G0XhVX56C5I5czFTSlRZEnGEDbpsFR9tP4OtG/eSLsr
L6bDRHin2HxVbolDF1BjfvmrbZsxo3o64JQ/n6n0fybdX+mERXIXkDj36SGuJNv0
Ynqb7CdRJAejG3QC5jvJRrP9GczYhmgr4s/MH/t8U7RYuDIRjHVPwKlOCBcNrr9J
CNTcUNxBqLqXHBvOPz/S655Mk/nxmzrl8QZlmQ9AAxqOxN+Kya5mBbQwl0xBhn1p
9Lffo0pKjpQpFP+kS0q3LAQIlvSCZTaNzSOC4o/u8aj8IfTmpykSRJAEXUBWN2ve
3YEXyJpiNL6dgrE60aYJRb5gCsd8ZMwWyYyykJS4ZX6nKB8xRboP1exR+iFBPmo2
4MPw2PiuPOnofnOHRjkvNO77TgniNQdPN0YPvsgNBvfh4g4yzxD5uErJFJTudywN
uZmMMCQFfTocONq9YTYLUerULpTYm0mMqTEW9eU9uMr4tJWOafeG+nzrlEtZzORN
Rdq0ofM4cx6rzm2fHvgQhnRrT4frlCCTfyWax2jJV7qTmhZhFX1/CQ/LCydM9J/n
wKkGbRRK2b6J5uGEPlt2auo0kspPkQnKYCNdOYTtTn0NzUCWtT0ht3f0006nuDVk
UaF87jl4VPa9d9ibYLaQSnEkyIHRohaaN7klxQrmHwWsigUAc2PjeogxoTP3zAjk
oToWQcTdtBQ0vYg23hfqkPbNBY7EzBVp5yHCmTWaCkY95dtwgYp/2wpCPjE9pyVH
52fiwRmLZNwcxzPjNKRpXVlNhsch9xYwDtDMXXrcb9iym+QJcS9/ZZYII/iVgh9x
nVI2uqg0t33YjE5U8HmllzYggAsSVcrsqg5NhItMq48K1oxy3JymkPsy9NLNFdpO
J6ckc002906r3mh6coBvTcAa263zCrXO0AOkVf4GtMlZNfHgH9UsN0byhpG3fS6B
3fEMZQXd5m+4DDUNdR3GUa5AcA7LrZhC4ke8SlUIWmoM2EZIc486XXGQ0rziKXPT
lulO2br1+Dk7ELCSpWjj50yJTBf1JFwMedeXIp6dkz0DJwVjPqlQoIfKcViI7rTP
/i6ym0p0VrtsTNwgs2La1iBcMCWgUk31XsZbyT5ApDYkrUv0QTbYD+6iuDkYPRUX
p1bfXO/bB5Lk3jsqq0qshCfcj+Is2SMoUiQRuL+zzGphCAdt2q68eiMneGjwqMIT
V1FnAzyHzVuOCDypDhy09jcz6I2OkE03iOrNQB4l419+PEqVv5JYxv1MEFgyWxEI
4irwE4V7zKE5a9Ubb9SpZx+zixxKAslri41L/QQkPXOAn5jcQtrqh8Oy+ZA5Zrbu
xEhJHOdGCcEkcqAudSWJ9H/a2UZBplXmmefBWNzIpufWnEuqVJjEnQz3CqRH50gN
nF2lceinZHxTbl2UVorT4bdDJdJiiqqYOjg9zSHU7/++lXgLimDH0GGNIp/3z/JN
u/mE4vC/sfOVYDeQPfZISO0t2EvHGaOygckFTVtt3a5wzpeFXCpJ8HEVIBbsVhaJ
5EEiLbMLUzyfT0emmfxl92bwCMbX8Y1OecBtDwp/ineh+JXFlm3rv9ujxYLCe3rb
7sJuhlXsjZa8hfyttqWZHTsNqRQjibg68Usn4I5OwyFd2wVh1kW+pbGQYPwPy24H
k5va1j6WAbFX46BbY0bIvVT5M6bZeoO415YbtQYRO3MTzlrFcg999NmWeFjT+v0R
mkfU7dv1vMQFy28H7j7id6ugiO4tCi1FkFowXhl/e0UxNYuYvJRZQV9qmlPBFfan
nMKuoQw3+IJMoWtudMM8ZNqKu/rd4v2eLVao6FDlh4n2Y+8xUo9S85xLQ3csD+tz
qfA0QKJS0zatlcBbBVzw+migTQeV+N+EllpFmB0D0U2YFfrYJJpNA2GK7y3jKGfE
d3V1zdjpNrL8AW+TFSa2F6rVKAks3ZXLsV/ksBVk2g7e/Q6JDCmyKbIf9jQ5g5hr
Pwax1h/M2leSzf8Ub/1a0Dxzf6CQdC4u67wlh03kgWotcIwH9Uw+lsoSIufmKrOt
+IStiDmlRn15kgV24LDDg4UKKRe40euRr7V3+seQeJOpFHtZFlf6HHvIC+kay3ZN
xJ+zANpyjABc6DyKHpxDv4zZjzn5eMSAiC1Q5+YSSzWc692m9Tic3eVhMl/HBVvh
f8rXDhRU5kEolrndnLa/OLAowAjXvPMSwNeVGgkNPuN3pglkjV6HNgKhaj1RjntR
M8JjbbzchKdG2yBfGszbAXIyGD//V2y5SlHXarLZsAoS0kYJvdny3DYuX1yDedF2
ChDlztcIcs+a7fG79t8Ld/7lux0kP8VaCuJ7ti2aHeCaliFsknIw+6+m79AChY7S
VCXP3dK2kwXPvhaSWwDVSSSLEosYfeh4JHmsEN1cpFLKTamBcVu4/zCUkXThWcmF
l5/gVXv5FYvBqW2xiWVRK342Nuj6MNTwi/pmj848EPwNxkntlgMjrmVHKSiGQBGp
4uCfA894Ybee0s/R/8j+wcwz2hCS0Xm5XLZ5kTb+pasy0qwOZqyVO0afEwMJpbbK
E3kGvpHJwjI5clvlNelqh30S88RmqNcyPSIu3iR6LF1VzPK6h8rdH/YTkwX2WwPf
I/3wBGIcH9GYZTGjuiERBr2nqlurzucLFbv72qDLN+v+pWpgSJB4FPLMsaLyYTiM
DcH/BxQT5z7VFGQJG6la7huBrKg89RQQvBOib8tIB5wSA2gPRgH9Tt4AX0UjI3gq
R3bx26pY6kT1rZyeRUPP1mnCNYiAcZpCB3/Gk3gh21A=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TsqgCAJG7npBGvirboIvVXD8DlqC23hgPJPUNKyoWA1XJyEhiOpifRehfUsFp6cF
mjOqHht43qnkj+//OySGCF9AASCautkedpMeZHJ931HFdO3keozk/arSLEQQFofL
P+fdL5ZI6EzaWEItBZ2/eCTh0q1dKkJOwYJA+8AmbT2bGFHYCk5t3kCwQOYqGEdu
IIA6IIeuGXNAUPMG+jMLO30YqRNQkdosnpZreLvRxeAVsvgiIkWN+jETkcQWQo0T
DEDFIxZYigrhi+HTd5y/T9oebXUep3rk+W2bFQZEtbv9FxkILEvl3yts8Ko743zG
Y+bmONsl0tofrurrgkc0+A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9504 )
`pragma protect data_block
rLMyZ6eDwCUr0PmV2l6bALajT5O8GkjmK1nEIX8eeH+j/+kbWQzq52P0rBVvjKCG
eL/C9WYdN4kgIf1IbSl4XWYkizm/PzieE5ByqXr2n3HIuUj4bt4edCJoZtTgrLkh
Acyf8AqRZP7uNA111raG+MvrRADyNXfnjl/OL/aElJCn6YkY5WXUzsKvihchc4aj
3CJSjq6kMJVl4bZYkcBvtDJb/oZZZ+HboIZoBpcik/1yJlpjRH9o0k701NNl+JDs
TCt9vTxsLe3UqNuzbYGA9WLCHo3Rv8abApO6f0pT98mHbfIzDDt0rSgkhQ4PGD2d
DRg7VmuVoLEclGOhxgCgx5JC5hgderHgXmYcb5BETvModYN6hqCg8GQAZuhcWtQO
hLnZqJdS71+bJirWoKeiqMo8O8VQ4zqTxQkJJHwZ8X4tsjTo4hFR3B41Er1SWrbr
Bx3YGzCT7mPzOPsmXZHQh6MW1fxX2Wu8puDTP9S0UdmHIrfINm7Du0pPJDAsQ8tK
zlISkLB9e/5tcJGYqTxGxI62TPja75cQCL2Qfj1+66O7OoE/rK7KDGwL5WwTjbYG
QIxlyMCKZMXXvuLAqgJ6sRWOh/rMsBQLQ2cd9+jH/SkyMYYKmNhqPeH0ZlLNHCDd
i9nkQbaGAsdbFsP7HX3kspw8sVcQld5Y21Fm95AssgQweCO13ywPoisjNPTlgy9e
3od2dDPT+EHjKfuBPwbUq+zKXPIer5414uzO0a9bV5zLTWq6IBgQKfrzceLG9sol
wNz62j14usoSOLkoON35qR+/Q7osI/dYTCsJxlePbwllPrzlQJSUwjXrn+Srf1vV
H34LpCvtIlhfTPqGiFFrEbJgWN3aAxj1ekGQezFseuSnWW9k+LM2YMYGqD5REbxd
rS3qaH9zlCUAAlpHU6/ZhuxWUHGKD8AcJ2pyb7SVG80qSIEpZIQagXFpSBesQNzr
1fhmepFl+L9shteHmx78DbVeVrTWjyTXsNQTZ7I1SgfhuCB8gqaZ+l/fSTAyHGRT
7gqzmAXQx8xGAsEFmkyyIIYTbIbjcTOsHTIEpR/aQaJd4ROeOaJgYg2EHG3b4i9z
fOGRQv3omTZX+K+8NcJOBCO8BUjWiosUwQatH6vVxwVyfvAQ1eSmplw642pYd8Fn
QkFTnLzpd6FDOGiFhQ4npEs+OPdJ27YphMmKh9miqYkdnftxZw4kYq6SrObzyUBa
Aq0kwmaQKtVfeyAEQhhnuTeleA937MXBFGF7jh4A+3PPNj5aCmlKgEnSC2/seyTP
3RpyLzq8KJKFA0FdaZ7yTZHdfC2HGbXQ4jgNZlkIJ9X29AUMQ1s56/5yfR1f8Jep
XVdc3faoTUu8ril3yg0wXPX7T6BIYAOv7qssPQrAbMVDk23WXbFL6M7tf8t6ifSr
UvO6idndgHehvFi6SOp+crqwxJ3EJDyB3BPDiAelE4i16cHf2B/l8rdMdgOUTgBt
PiyHw6OTDc4Ox99n6jSeImFQO1n0wZNjTw+gDLajlbq6+xI8BU4YwTFPhXpFyWxM
iXQkmjRDMl/f7ap2gRGsmWm84jDUOyxIy4qcfxEcJyquYuxTO72GBMYDt3LvY0PR
O8jNueyqD7cxTipW6o88M5MKpWdmRkLN9WRirU234eLmthE6zj5m1FL8+p3do/XW
dFz1maDqhw5J3KQ/z+QotbVOD3LTUT4oYriFuKT+9Pj/7sNuUO1Vb8WDwjeRUH3d
oz1+wXBNUVw1cUEQ2CNZz2GDFxegToZCNjFA1hc3T4eDfVBjn/4ptZ6fGW1bhcuQ
ImHgZrXjCQAeARRxvb1dWnlfNOR4Af/RjRk/sDoGnkHTZEGXKbtwIvqSuHQ9v9SI
DsU5VYsx3ZeTaLdA9XI3rM4yqfmymiFr6HhIBzrlq6cVyUowLwzh3YI2nSwwp1OU
oORJlo7i1IPNTDJo4/BhQlLZTsD328V5D+nECbqiweXD7jYTbikjc0JrQTUSV0A2
2+zwuNaD/RY/LzUGRrp4bKIPUU5OUrsf8Tu1t+CYDdJC4qO7Y9kKXLEMgskNtVv8
ijL4ORDxnF5K7xJrnrVoAVJAXOC/09emgEj/tNFgOwHcpUQdjkpJOJDuLPISqB82
9iMP8Qp8d3nSL/XrbXeDQvVdkbGV067hvjxArpLjuJ0sNcHPktLj8M0hFOJsI/TS
wYIh0YfBuHlQdCh2LZ7co+PVKggWOlMFRSnyXNszVIeTR6kxqhaMPF7P368OCKH6
oBlkW3Nt/fZhe0Vq5ihKcglIXRu3Bia+w9SlVOwHo8avSoGXG8iXxqlwM1TMOnIP
8/TvQKwTLSdFMgC4NgywuIsvcjoKpByPji5AqiYaz9IyqvRml8TBKCDXALLL3l5s
Fdc3l5AzlPpwDWSupCpLFcKmQcIZZHRso/nlB+UItqEPXh7fhYHmzCGXxUed7c3e
ouqS0yCnV26yfNWQkuoZkAgKx+bAM+Wp2VxbZiq9uxhcl5Nle6GLIPvrvT/kZPAd
cZApIHGKtyQCRUotmQZtAfwxGXeYwpL575E7rteEBCV0XdRQF1McEMxYx9mer0QO
Q0jxqS59JqHpVVJav7sEh1TWTgUQYGejwZP36x8NEOEE32YVZztUqqie4TzLeRvI
FL8pAmpHvSvMeIQMsPUwOHQEhqLXA/qqZEX4aK2qZwXzhZBwzj22/mdetQ/rNc3m
0H08GSB0ON77fKeMtZLu7N1FMyXkF5LcLdEH7u4l9nCjDiLanUsz+tTnJT0DZKPl
O852kDg1ig78jGhbVkxomFdjFEKE0IfcnycfYLNdWs1/Ao04jHO7kzyM05G806zl
+QJVNgGPc5mm4AKfBNAcOsMWgwWF9pgdRJj0p4spxiP5QeK9eakyNAoc4dkBrJFN
jJghQNWsusMYsX8TwNLHNo29xW8G6NyvaUXnWIGzvcSf1rZY4nd45aikQ6n+4Cd+
Qa4N43Q5xkcO8b++jsGlnPF5VwsfMM0OFk2kYhj/RxLBSGsS7UlT28Qz2rFdwHhK
Y3CmneLx75bsH9kUXUndGohI2rbFhg+kceJLvCYS9Iq8cwPIBdlWvhei8/0iol3b
Htg2BAv8UW6IgDQHBUlitVM/vLURtDBIcIlZxnbClQVLoAuPNcoEE1PBQKauog56
PFE42MeqCI/6xCl8MS2tW3ogt+aTE9xKPwiPQKQ+zZ/7LnDBmd1ZLDW4ziUhJm88
R9NB/nk/sYfYzaOO/lwSp/lznYVuqkS6ufsfNb8nvGbg40mXfLhnPCyW9dt2dAO6
mitekD1iEsYkypzaH7Ao9wHQmCNMEGu7v4m2WGuvFqs84hCfz3EqL68tIYQmtqj/
mhcATV+3Obc+tbeGXL0GAu7TS732i+uPhlgX0/YhAo2Zn3R3NKMfnSMQ5QhqGxZs
xk8oIGl+vVCCuJw8O4niaDsvfbxdnkECh4HnLcW3DWqVl8cM0NgvlGKSiR1WgtZa
bZrCetkOf8CpWd2ovAF9SA7FwifTICprR7rGH7zm9xHZ/T8UWKzJcQUK1x6zNJzq
8dm9qUjJAM4kRUS2hQJGG/nr+d+lXffznVfnVWnpiv0PlhinTZ4MF+QdZ9lnVLkx
AbIJr80vzhC6X95/oogzw8RRLBmCxRMG+ymvBkeI35F9dsGrm2S6wGDu/XdeynoU
7vl6qSBSkmnO6oOIsTwmIdwWA0mfpL7JiERlhSyCd6W1NSytZoxjA08r751TT3BU
/UzQcgw/sY78qkkxpeRjKuN41ynILATlVMErto5dq5ZumpxPCu2kxc8WnKMJx4sm
3c3/eaX9KCv4Fg35uXzxsq/YZpqYdnzqK6uBpA5nKn6FYwFoavNKCKmPfneoCdSa
7qQIq1JgwEr3iABANKCXrfPLdhC1tWwWBdNw9FPpa21KmYNsgIGKdInjNzYPFLtJ
e4NXGEh4PDdGFCt5UOizS5qlzzyTMGoWQ37tfxCHSQtM+QmBVEAYg4MB8uuzm9X+
ttnw2q7QvZWYmaRUmYe/lU44jgULYpNLIoW75x6/ALdMrlc1s0Oqow1eNWmcbcWf
77qUqNeuV8T16OE8TW8rKN6JorcXP0U7XNZQRdDqRhZ0mEODgk0cBa7lW5DmkJEN
Qm571ovpGgEBxkeVnda/hkfsGZU2px+NI9ZJDPNUrkoSh8GAvZpEp7ZQkBAeA+tu
zQphW+/dE+rQNjTNCNcatsmC8630f2YhFvIylK6ryce+u5VRZCuKfYq8JWNoUGw4
QlX/BTxFVGq1cQ0KL5jydKzHuhdV6UlJAnAFQopLM8PsFyWQkCSiGNrvBz6/WBS7
OeQ+galKP7an4+CwvkOOb1kUlQedPYy+CFtppf39RpUZZBChbrItK3JsBqgDuC3W
X0Os1+U4yJXLcQRyVbsCR/Z1aWRiC2A/YjpBJ8MwK0dHB4sSEyp4M9p8HzntdStG
enln9T+l9uCkgfE0C3ATuMuEtn4DIFFlXXKZYIFYuVOHSnK+OsZeEWXoQUmstuc/
i5RiMXt1IF3qk2o4Hnp7r1I6T6ODr3rL0acfBq7hlcJ3HG6a7UbKzpIkswJh8IOo
tikNekYt3fhniuIiVrRe1A7cGo6wiePhEwAGAb2zzPZ9kr7YDbFtpjP5aRArfi5w
lkLljWhdi0V9QcR6c7SlCFUMquVY+Z6Mk+KhU/ynB2uS7h2J8frI6Vfj20tNAGCi
z9ipvoMB6CV4jqGrQqILpBjc8iKwLGyvsRN8+CvaD3iu0WkkqbO7LUQ6aZ1PIlzn
u67JlGB9DEex7F4EicG1maGWCM5WDG//fyrhM2jHxut0P693+zBYNV/wO04wSBGU
Qni++3EaSfxi2o+F8MIdqoibHVHj78Upiylzxzqr9eVgGvmOxfPhwaGiHRMba19j
xRK74jBC/odBQWC9i1DHHEEEyrMQtJXN43qZF6NOUFxN3Oh+N/HjCQS1FxQ/NFap
UAdKDQZm65IEzJQbNACv5+MLJrqPbELcIFXYdPJKJbYUYErX2M6yfQysXqIlCSmr
zSPtFejFl2GqQQHFJ209n6eWHKQy9OBQ1CTsxqqWdILAxmbgg1462c5agITEUlwP
PVxSiNmIXez3K7hYdai6QNkAt2ZgCW2Yk1y5/yBZ7w0DoEcj/507yUyFj6Sdzi09
l0s85wlEc8qFlFGquy4NTnDkJ+Cq7Lsfw2kmnLUN9sZ3JMqc6ebKUBtPawXsef4g
o2D7T6znuaXSIRni13yTxR8Yx58S8+SI4HkC58fibwQGlgXxpjoWEH6QF3L8aInX
rCwC6oMhXw2QdnhY0ijLHTwZNxB0fO02mFpDHpVEwy8qr3iDj0rtwcDtEi+8NNM/
s+97rb1ngRJBJHNm++oFdzk91NSzBtI/Co/VpnAJEll8Xu6GLmvwZlhlfXBodUi4
npsDz+hAoo24ilY2T/k90fi8Cmpm9nCLyK5wpR9iMT+Zc3vMqIYtK7Mbbk4bzPCc
4dVDjt9SC52BztAH8o7EcTJEuEI/0Z03wqG11mf5gj61tQmeEN0m/3siH6vnSnHZ
QkJDcldceWD6zu4hxKwVmcevtYJbZz3orRPh5bNo8qXPtVbMimGciO/wFyaTBeiV
njsKdp2CCYPNszUI/YdTedohKiTTm3vrXSDg9oLK1ilrRimwxotFZvHltlDjg++6
gFqfcnWLE3itQ3BFUiyWA3NOdsPpJFrJq/sUXuX2qW1c7Il0+aPbZFJdMFAmCvno
8SofxJ0fblxqh/toI36K9R3bbEcn+V4YhGS+y93zwIeZVSzzpmyu+t26q+eVCMGb
oDAtG1BS0DtcuKcBPSu1uGIuKaQrd+xnIZrKveVHe3xsY/WnMGllO1DdAD4Czm7D
MssDTX8oZFTqSxeGAkNlU28N9msuQ6bDfJWzt0DFohZ2K/4zL7Dh6yLmFMJBJepx
RmIhkvecI16NbmGxbU72ENOiSgu2o8YdcczjMdWnYFOZifmtj+fADey7EwkAork4
bKfP5h4xQjs5UcU9tsZsHPhn9uKYsBQjqJpJJmPboGxusZ5zbk4SRdFwQIDeMX3u
BZJJ8miSx9nrAVJg7J5vZ4Vdy+hedV9d1EXCQP9sokk6xN2v+FdyMfNZ8WBQPzNK
kEXcFEV4jmr1DvyrPezARwprg8akEDAAFLAhIej8xR/oXRNv9lYYnud/cJ3kQfOk
IcrZz1ko9owi4SvT/yTk0tIo35KvUEaNt0VIULlIo9fz4bkhM/WPoEGVErqjILtw
10RxRJgxFfa/r4TilJl6wyHSn+wbmF5PbOAq/W/Dle708ze+qPn73bX7dnLdSelr
NO96TiKeUMVZhJDfGi7sEMhnjLHhkC6ZMPyhbomQ5CSCSHEY0P11N794I5A96TQ5
nxzAn7FLmBxQwSXzBnaOCS0wEFAB3wVnM6sSj/DAhvhW0C7MJwaZa1wKUCLAqJcF
SjtVpzH8hVyqWaMsSesEd7giQHnyZlFhemWtXk7AGjG/YXItuUyp1j1/2SoDtJXl
0kYZ+f0FtVWmRsbsRCwWeOGT6+APKfgPgvrOFfvbK3uzn8tMODG1b6az4oNOVgS2
g9p8KjcfzNjLZQq1xSU564R6bcoNM2GISuZawrXvBGQmbQUIj4S8KDoKNndgi/dh
Pd5PqYfvxqZjFJdrgMwD/88qMBTl0ZPVMYv5sFjc8Ylq6sqQmCjv2BqoOd5e3vYd
GB+V+CbIBo3QS0NuOZn46H7+pV4vOrdXm/EBSU3Sz9k00tSU+EBe3O2zFIyVmfIP
mDt/kk2i4dSEUk2BOlqBgiolrXUvrnxVkR/Ms0QDRLSZdAGhP2drfirzNiIcwinr
PDCM5jSCJ+CJwtpWj1yha+zhU2M64k66hpe64W6zG1DTXGEEvLn3pTlgxuJdK/xV
YOtoD0G4qSSEEE/sEZEEXU6umkyl4u2t03SisaYzDJVsmC9AFN+g4bJyi97zCZ/0
UQ6KaBz1vARUI2vhWYwMEMFxluj0Y91fWFQqsQZA6x/G6i/apuI0WHYO0mYbqmuW
vX+EUx3vNg1/ps83RPj1366dI0mzyEaq0Ukvc8e5MOZmY+9xxMqHDyuF8Zw36Pv1
rtB3XjysXBiItZxBp3KcnewgSHXUIV4Jcu0OVDfztPA1dfhPN/vujGYH7lqei2qu
kXhaPxEqi8zcc5iUTo3AgKXbIARkIin9u3xxlZDrxhP2JaQXIa19O2NDCyNh8clu
khVMjCxkiI+L0OUVr91JFmP5xPRD3/Dw98+DJxFlcxbZpo6AfKQKVH+/l7k5U1Um
9aKDNYRopenbeRRLe7pE5elo+3ff/+38SzbmomnigA525dvQM59fDuaKDr2Lf5ZI
lcm9l3J3zGkojVdcSyPa8yC039nc4v9zX47DEQ7Si8yJVYxW8UZI9/PdV2kk3j8n
rcGlAKlK2GJ2tKyrLwWO1Rd6+Zs5UkJLj30gXqQcLrig6Vtxy7uVoiI9khdmCURm
UiFdjquHeof+dxJqhQvkdgFxMCZzqYJ2Jsi5p8tu5ahQnyO7nLZS84zbjaukzhY9
tUrneTw9jjMba1mClONEp6nux/CtjgnE82D6/8WDkblfaDSILR0IBmV9P+0Nv/GW
ZXsTGC31IMX4UsEcSrofvs0n//N59uOOy/OVDehvq0McSDcv4DmBlA1B01pcCRr0
rFs7k7rujxfgZFEQ8iu3s3wzFRg189f6qXMl42oTsDEq8ETawOOBzICprcbEXv8g
EIXiKQ/K+Af9PZ8COMpfJW7A692XKn2D16XfHwm4LOPBEdopcZREa2sQ3lNtXOQ1
Uv/XZNGBES3PstLnFaG2e3Hti4XlfJAQ5cHt/+0i/C5jY2/HI5kYbJ/WV5miXiTf
LPr7Tkd2os47dcssG6m7qiuPi80MtMeyjnzdgsJCRC484IjPrBhtaz6DmIlV+c8o
5GH9IdwQ6dNJpYNgGipwqH/Ir9RVZSxVJ/qb1AunVurCpw5c5jMvJ/Ny4VHJPr0b
xpn2mc4qI0Xpens0fCUmW0c/Fd4KBQZKZrnLRHVzFlYX/+mCtrFX3v+YSUJj9rXB
Vw9JxuQDoOUl5E0pVbKXwX8PNkhfFO+je2tQZaWzawRWp+Qe3Zd7b3OkAYGMNcuL
ylQBW6xr8BX9nQHqVrnRsZpkxFUdnK9PY/afYuOtfsqN5C8hizA3mWdIEdeIcJtw
Xp/QpbLBcsp8TzO/EAc06QmRyrSnKmqz0GsvLWyqh31/2gu46L19GQxF9i4My9gb
Z/KPa5eCdTrG/jCc+SDjF8KBRcebov+KJMx/W3eaZRpxA/9eVyxZMaqhNmVrWgxR
uskTp1Y8cyG0cWYGgPFDV+FmI4rOhZgFx1oufUxu4fWG672JawMvD945Ae8invfs
m0L5NWCEZXiizyKoiYOz/HYfpZe+rguORKybCv631whWJ579nPLW4qDiEDpyN8S5
uVYZg3fczKV397ge1MFnNfqMGRHGG40131L5/AUmwYLlA5LhCYus9doNTAEbdg+o
Pbf+DEOZLdzkCfVWPoYTCS5P+4vPS5QuhL6wn0GYE6GAj3yyAyWRy1GmsMZLUMmg
DXNwi/dzsipEmJgD+TmIFdSNDMsexG0AcS2ccGbMCppsgyPG8quIenQNwsw3G3T+
qYGAqxZrL0rNHOypkoPAAeqCuxTgpl5VrNESMTRGG9iMwQYbxD9rK08pOGpIGNkb
5yH7CpTO9cIQ9Lwd2d8OeD1kN7Fq2Hmu/tJt4ZRt94KraK3YVHuzXyZ991VFlzLJ
yg6CqeBhGkt+5jkLW3GHkK6kmLYu0igtAghLIji4Lr9xi6+T1BrwPN6XCYnb8AxQ
Jf3v7Z0IIx/Uqp+Y1e8m797VkPskNh/e/9XLoVtY7u00OwVWGsiNjrXMM7wIpXjq
4GgBXc6KgHdQvQd9/ebXNv4p7y0DUwVQ2KILoKjIxTaqOVIebQMXZpKQZ4mkDZZN
nrCpL+3AqoI1BAki7TqteK6FZ5Bjru4jIxE+l44aDpVzAjiP2jZEY0EC9S70f2OU
M6vy4jAJAgFfiKtc756rZdrmBpgdgKknOCTwmIgDY/d6OJbZEwoIyyLT7AlZLxrN
gCC9G60IRRP7Lj/1UwzAAiC9+fLuyrFTu1EU8F8Arqty0k4GQ3w1Lzcf22zBSJAm
8FcN9z/X9YUJYA+VIheAoauCrYasm6X3PZ2z6TjTwBgwe+HyDVT5+fmdV929oSgK
JzsY44fQTu1hRx4g2w/tPkIA6YR/q7vZr/mjLxbRuvQxJtjNe5ym/GR0Q960apd7
4ZYqguwNvceDDk5Z3uyIv2o5KEqYAsPpzbKMcTIY4TQkAOnTBlVRVSbQmwd/fuZe
3/3JBDSGmqttdJA+wcsyfNt79QQZOsLUAQWfQN5iRYj2qUwJWaHqdcCB0PUDsEMj
mWhaRC7TTlxnkeV4djD/KCahgvvH6upd1sdCzzu0DyB4bCz8EWvm/xhKRA1LlJhP
SQd9WiL8xXAd1Kyia5aW2frMwYK5KcuVnxDvfh1v/JiKTy27hA08eEdsnZPaWblr
c+GmGd/2EwW9yYXsLlZC4B9itoimNoyJR+j7cXvzxBq/aV/kdEKxlosg/lL6N5aY
Q5QbsQ4BAxDPXCPEoNNY0iTBhl3+aiuAA2YAirTdZ5cRQstqlVUqU1WUlaqTY/Xr
dXKL7n8C8ebvcxpPuHgiBPl53IzKuNmv2kLae8niAtpzNVWKP9UQEbexBHp/XJQD
hbq3fI/dnuFp3RwgoqBf7EL0C1z8n6KR103P2F+tj5zgpCU1lpou7KU/ViF+nwTH
a7RQqcXWH1IrZPYuw65qHacnCG1l33ouDv8U8QgEyurQRpA0K/x+qvCt2kmABAL/
TS6jNYlmTYIAy4X5FuTApZl7XUjdCYHOYkUxtv42jaXuONoN4jZvw40EkGG/RDHa
mhFHFrjSM2t9Nj4bGVa2rYebYZj80pyPlyFCsljSKJKEFtGWZIpkbaYMfPTbaaws
OSpzx2guHmVr5j4WQ/exd37PoKL0jeNek3pAiruYhswqgKRqNF+Ep1i7FV0rUNAM
CQOmc2il+ceSPtgrZ8Olj91vl/kDLauMukb54Hfg2fCqk8GfSrTokjgbZa9tGxrU
FpGKpFyYwO8u9NjDGrsIgDS7AmM6lDLJGBm4B05t1yYes6OabKx8L4OzRf+jZZnQ
NEbCAzsSuzPk9b+269OqFa8tCPIJ+YLvhv/SJIowUTHt5Bqbiptqh6OzquR98z45
5WytYGw3VVsTf7LJtUY9Xif/tMvrVIFtkDXb3kRCySB0u9WEs2gsJZryJEBVXev7
dCKFhlc6VZrK/o708rrF5Iss3tBluFyxK0gXEOkcgrU5EYazYPfzK4eUj1Qi1Y53
FAVdJve6IDaiZCbcJyHffVvjmBzaA1PR0zTwaEJmHI1/2CuzZtiRdYEpdRH7ABZd
0DGGNjJDJYU0FBvv/ARBNoEfWToMA9evtUDhhJrJoaBvwzHaynCi6fEDqXE4hFM+
6sL+bsxgBTy+U09Jprr8UaOCCVHYbz80qrXkNcX2Q2rt/0PI7Ape2KhW3DYG1xR5
TnwcsUOp2WOINKgDv9epSdQlBE9fYlLzBPiRf1s9rgC4bZ5ICtoU6sqPmkzayXht
hYW1z61lAR6EOh2+CDe20f+X0QmJEdhB+3PAmQbLndZd5cF41K8kXJWw43AouJ5l
/+SaTGjIZL7p+RVPmQwg4+6rQtll9LA1zGDt5OzG17o2AV7XN5WH+ZKiClfWBuiQ
v5XwnwbAuArDbUZcuoAYU/DoZGb+eTZa+XWa8G99qyrJ7Jnqz1mZREhdcxJWuj2w
VKXi9WwRFlYf7c03rg6emLzGB/dYpnbWFmsAUc9mwRK3x3vEJ02TUCGv9g234p4W
ioteUdFzCQZ1wzj23vgbHxh9+PMwPhRr7H/SKRxkDYSK/6my+ng4T468CdebhwnA
GZEIUwgEEBwcZBlJmrMRFuiRTFfg4BaqpM6P9I4rkwfDURDM36ykgMpIwlnZR7UV
hMRhoUD9UwkiTIBf0jjBTVc0xizRC9aA2+kLw1SR6Kx9BgUI3C3YCqPcwD8uDWGm
kZIabw4wPQyV22YraqnZB3+NeKe15X3SE8pfs+W75Hz+Y25WDOm+9KPFj5ubB55U
F+g46Qn3dPaiKgu2y2BIM95zh3P3tK3A2kotyOr+tjXYaTAUHxpj1Kj82u7mTH0W
6xVm6c02qOsr55IgWMhGjlgF2ys8D7RrYUXP8EPPYqH8EqC2ea4xbd7qVQ9dqDCb
hUWeGYkBoctQqNFdNuisnaE05YXNOkKUgmsDEqioolB5JBMRGW7SO26tDe/C4bn+
ryVdMc+I66gJ4SXBvRe+C/3SsN20WOOtwIdUp2IDGk4ckJiZ0IPuZhSzAqamhbJ+
y+ImJ23AXrwJmZlNW9RdFb3GuyDcn31KOtVuVDdTf8Tg9dcrP1Zn02DjiPFI9GSQ
NCaBZPdh4NeJ1vHW1WiSP7pdWaspKzAvPN2qTd8JQF6bz3j6E93qcu1nRgkUDNis
PzVQ9jWVuy6yrVEOXHsB+ZrrF56Udci7NbLH1pNgLCIo0flqIeI3/MHXuxw0YAwV
0VEhrfTPhy3CITo3b9cfVArnN0L3PQuICcRqvepYKsvLl5k/HHHtX85uhEUZIXW5
nkxCzq2V+yOltUn2lNXeHvdFUx48CZBKWlrPkJ3Go66cWJ0XMfMzM2X5yaDTcTAY
738ZLKJy15Jfy02uels4K0irIMlCpQ94NltTaQFngnhmarM2yLXqsy0+E9Onhvne
mS31uY/2KBEh63UKpg0GvG+2K585wZkbKUn7PX61SX8lkg9abvSoLYxUcri7/9n/
2mpGR/I2tWMO+5dlIy4P5AaPNHGsSketoJtP5sqXat73l0JajfGy95XvBEHHg6Q5
PNg6PCzyO5/IQEF1LD64gPnIo7LI1uTJeobj5TZONweJW5KTLAh2xvu9fZm6XCbH
+DaRya7hGOoBf075CCOvYbKAm/BOnCKL+YysyDF5l0iwFQ4eF3v4O48EmbB4MblL
c4JSOV1biHtmh4i+1fCwJ0uBbVkl/GNe35742IY+j+kcieZCrsgpOeO+kaM55j8y
yEl43q6wefD/jgRMUeXtEYPzr5OKDFQ18oeF9h6mAktNK/HxP85MBDzCj3V7laW+
HteOonYZ72J69C/V0Nanpm6Ki0f13TvxmIl+iNhN8pEgOGth9/QTYvs71wpsHfMN
fOTj4rgiE03sYeEzF1jNcKpL0Ydukt3Ts+TVQKB77vkQx2drMnnr/TF7RDfzNteH
h2nTyFI0kIcnt9UXyrYx4BrumD9uh8H2kRMtcKqAejcpz1Fu2ZwWMu3shFLre2QV
xBI5wm3mQAAyAtWhmD/7bmjJ0uRss/wcJA/OhFFKa9zQMz3j2+dW73XP/PUND8Hk
Ga+ZYHV2Cy5jnJCraOTxzD+pB2I7n9guZ4X3VDipovtq2N05oJuM5AG5ot53aqRQ
VaqMw5XHKhKoa6XNoKr7bIeiNhTZDb7eD32aqg557KBXfjw/vjIqudYksc/HzKZ1
XtvIs6o3nCvsUQW3AieQLXqZx5rs+mfTGpZ6WqWwL4lRzIEaxnK9bJukJWNegxdq
oHvUkVV4w/e3H5WE9aJ8gpSv+rcY6lo71P1HVZLszzv11zV2dsZ/NO8s1aWIhLbQ
gJ0OwMRoxKytkG1wXNDR1afdnrLLeWyb5BeUA3bJWXNqXV9JSgk/c31MCQraC6Wg
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ayrD9S1ZeURPmSWtRI6UZ5wp61UBaQ1IEmyMhAE5HFNg+Nw08Wo1gmSjDSmmRH7L
Im/di2VngNSeZ41jqsEYSjbug8CPrxgxQxs2OWn5nnz/OnPDKXHIELG/bOjqN9D6
o+EhGSdQWG/np1OIBrxbBQZHAzHrOtb+dCjncBQ6/4RuTAcZ4uZf5RVY7ohWnH6s
qt3iSNzyRa739c4u7uwJgQfhoxJM2k2BeKDuGvtdML/RCOLHuzvA/YZkSBjlr2S/
iINzgZXJE5007njB9ND1Kw8PP2sEHoLGT5QSa83XgggKAhojy2RDNwcFnJdT6Kwu
GujXpHAKKK3G3+l3nXfM4Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 944 )
`pragma protect data_block
WutshUV3EZqT7K+y8VxIiAlBmT+zfqtwz8LAi3Tt6wLvJkgQusHUz/r5Tu3iugGr
gQHchhYwwK0glNEQ2vgVLH50gTV/ZWhazMJC7+LERjVB7ezp9GlftqNfEyyfXw5c
yLO+r/3UXTDnGmFwaJItbrGl7b9uqFCuggLivmxaTFrWkt73sq1OyM+NrIC1eCJY
QL7b/ALMeLclLs3RB8fIfWSVcPxMBFL2YDPQaljesJQ0iiLklp8dtEClpZddkWSE
WNKwnBPWHUxwZreJmKIUKnLayEfj9vWLuX9yIrJKPgXNNUxfpyfNVY06PA3fQhuF
nXz9zJ4bApqw5VmBf7wBWoOefLqItnpxZOF4RVJXZRX9osdiIRmXl0PPBTXyE58z
LpWmWYCJ9ldSDQbwkUUapn4XxeyhOkdxrnrN9jcK0py6EwHc0IgvH9ZVXo8qYPui
iKrJavPyrjj9asY1rLxYBSUs9CP3e+OB0oeT4W9ytYXjPD/oOGI32dqltYBnMoOv
mhdCD+/t3ZphNBFGOSA34HPkA2XVr65h9CIPX/EO6h+H22vVCfh/II+70xtO9JOU
B7tx0nNmF5ETlq9rVDb0HxAmBjOKVTo/Z6E1KUZ3JTPjWywJQSdMxWJpEGWVfrpV
eJRjXU8vAFN/VvxNnAPQ1C4I8F7OBiqaXyX/8ne+KnplqrmfMl7TyW6fFhDm6Cny
Vg5kRhtRuqb7/lug2BVK8NyDWXEIhBuCKEnuO91iesLExWk6ceOEz+XIi32PUQme
k4WSnDlW+v+lzbpsR17QFqoh0pmr61oTphoeXkKaKMasJaXj8+eL+DuEkqCW5l3r
oENHc8jcG3Qz8BQf7hIOMwz9TKaPTZiZM98m/TFcnP+788yEijT8xTM2C8vXyfhG
brqZhiOqD15VKtKYt6Q3EEpjUX9ubHhH+us/JAkyhdzg7xDOfpH2hDPmNYoZcG1s
2TvRLWYoGrqeA6hR74nbv+glvhr6QssY8zW12wRvCmudSUpnl8PxXyAU8yaEK2l1
DbD97G3deUyhIUm18WRLTNP3Pu16vhY/T/ger+2UXX0nUDr/slv6Hm1G53ntgY+V
81k8Y25UlTo5LbemN94I+LAwcYOp8ylZYsq9e/VGf4UtkWgZ+yxXwOXfrL64kvhj
RZc8QzJFtlRQOs0BdCQc2b47lnR0p1B9Ri1X7QvIvFNbqPr7oFPL2lmqVXTeiLQ/
uflwDgsWPA2ig5KTqpuf4PBFMMJ7nsHTLY0XFRiLC9U=
`pragma protect end_protected

//pragma protect end
`undef IP_UUID
`undef IP_NAME_CONCAT
`undef IP_MODULE_NAME
